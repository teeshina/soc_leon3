library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;

library techmap;
use techmap.gencomp.all;


package gnssmem is

  type ram_type is array (0 to 65535) of std_logic_vector(7 downto 0);

  constant ram00 : ram_type;
  constant ram01 : ram_type;
  constant ram02 : ram_type;
  constant ram03 : ram_type;

  component InitRam is 
    port ( clk : in std_logic;
           ena : in std_logic_vector(3 downto 0);
           we : in std_logic_vector(3 downto 0);
           addr : in std_logic_vector(15 downto 0);
           di : in std_logic_vector(31 downto 0);
           do : out std_logic_vector(31 downto 0) );
  end component;

end;
package body gnssmem is

constant ram00 : ram_type := (
  X"00",  X"27",  X"10",  X"00",  X"00",  X"00",  X"B8",  X"01",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"25",  X"4C",  X"00",  X"00",  X"25",  X"50",  X"00",
  X"00",  X"25",  X"BC",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"98",  X"09",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"01",  X"00",  X"DC",  X"00",
  X"02",  X"00",  X"D8",  X"00",  X"03",  X"00",  X"D4",  X"00",
  X"04",  X"00",  X"D0",  X"00",  X"05",  X"00",  X"CC",  X"00",
  X"06",  X"00",  X"C8",  X"00",  X"07",  X"00",  X"C4",  X"00",
  X"08",  X"00",  X"C0",  X"00",  X"09",  X"00",  X"BC",  X"00",
  X"0A",  X"00",  X"B8",  X"00",  X"0B",  X"00",  X"B4",  X"00",
  X"0C",  X"00",  X"B0",  X"00",  X"0D",  X"00",  X"AC",  X"00",
  X"0E",  X"00",  X"A8",  X"00",  X"0F",  X"00",  X"A4",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"25",  X"90",  X"00",  X"00",  X"3B",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"25",  X"74",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"C0",  X"30",  X"60",  X"32",  X"98",  X"00",  X"02",  X"08",
  X"FF",  X"03",  X"32",  X"98",  X"00",  X"0F",  X"00",  X"0F",
  X"00",  X"C1",  X"00",  X"2D",  X"C4",  X"CF",  X"00",  X"93",
  X"00",  X"BE",  X"00",  X"EC",  X"00",  X"08",  X"00",  X"A0",
  X"30",  X"60",  X"00",  X"22",  X"30",  X"64",  X"2C",  X"2C",
  X"B4",  X"B8",  X"13",  X"02",  X"FF",  X"12",  X"0E",  X"00",
  X"64",  X"01",  X"02",  X"00",  X"02",  X"00",  X"00",  X"00",
  X"12",  X"F9",  X"01",  X"00",  X"00",  X"00",  X"06",  X"01",
  X"29",  X"BF",  X"60",  X"01",  X"60",  X"08",  X"00",  X"A0",
  X"08",  X"00",  X"A0",  X"00",  X"00",  X"00",  X"08",  X"32",
  X"29",  X"30",  X"60",  X"AD",  X"68",  X"32",  X"98",  X"00",
  X"09",  X"98",  X"00",  X"00",  X"00",  X"04",  X"00",  X"00",
  X"00",  X"08",  X"00",  X"A0",  X"08",  X"00",  X"08",  X"00",
  X"98",  X"48",  X"4C",  X"50",  X"54",  X"58",  X"44",  X"FC",
  X"48",  X"F8",  X"F8",  X"30",  X"80",  X"44",  X"01",  X"89",
  X"00",  X"08",  X"FC",  X"30",  X"8C",  X"30",  X"80",  X"FC",
  X"54",  X"00",  X"FC",  X"01",  X"00",  X"08",  X"00",  X"A0",
  X"30",  X"8C",  X"05",  X"00",  X"00",  X"08",  X"00",  X"A0",
  X"44",  X"44",  X"08",  X"00",  X"32",  X"00",  X"44",  X"00",
  X"44",  X"00",  X"08",  X"EF",  X"FF",  X"02",  X"08",  X"32",
  X"00",  X"44",  X"00",  X"44",  X"04",  X"44",  X"08",  X"02",
  X"02",  X"00",  X"18",  X"18",  X"00",  X"44",  X"08",  X"FF",
  X"44",  X"08",  X"44",  X"08",  X"00",  X"01",  X"FF",  X"FF",
  X"00",  X"0D",  X"00",  X"44",  X"00",  X"44",  X"00",  X"08",
  X"EF",  X"FF",  X"02",  X"08",  X"0D",  X"00",  X"44",  X"00",
  X"04",  X"00",  X"00",  X"01",  X"FF",  X"FF",  X"00",  X"D2",
  X"00",  X"00",  X"08",  X"00",  X"98",  X"44",  X"48",  X"4C",
  X"48",  X"F8",  X"44",  X"08",  X"4C",  X"01",  X"44",  X"08",
  X"44",  X"08",  X"00",  X"05",  X"00",  X"44",  X"00",  X"08",
  X"FC",  X"24",  X"00",  X"44",  X"04",  X"44",  X"04",  X"00",
  X"FC",  X"48",  X"03",  X"00",  X"00",  X"00",  X"00",  X"44",
  X"04",  X"01",  X"44",  X"04",  X"44",  X"04",  X"44",  X"04",
  X"01",  X"FF",  X"FF",  X"00",  X"06",  X"00",  X"44",  X"04",
  X"44",  X"04",  X"FC",  X"01",  X"FC",  X"01",  X"FC",  X"4C",
  X"02",  X"03",  X"00",  X"00",  X"FF",  X"00",  X"D5",  X"00",
  X"44",  X"08",  X"00",  X"0B",  X"00",  X"44",  X"00",  X"44",
  X"00",  X"08",  X"02",  X"10",  X"02",  X"08",  X"44",  X"68",
  X"00",  X"00",  X"08",  X"00",  X"A0",  X"44",  X"44",  X"00",
  X"00",  X"00",  X"44",  X"00",  X"47",  X"0C",  X"44",  X"04",
  X"44",  X"04",  X"44",  X"08",  X"44",  X"00",  X"10",  X"02",
  X"08",  X"00",  X"08",  X"00",  X"98",  X"44",  X"44",  X"00",
  X"00",  X"00",  X"44",  X"00",  X"42",  X"04",  X"44",  X"00",
  X"42",  X"00",  X"FC",  X"0B",  X"00",  X"44",  X"00",  X"FC",
  X"04",  X"01",  X"18",  X"FC",  X"01",  X"FC",  X"01",  X"FC",
  X"01",  X"03",  X"00",  X"00",  X"FF",  X"00",  X"EF",  X"00",
  X"44",  X"00",  X"D0",  X"40",  X"14",  X"44",  X"00",  X"0F",
  X"18",  X"00",  X"08",  X"00",  X"A0",  X"30",  X"80",  X"00",
  X"01",  X"30",  X"80",  X"00",  X"30",  X"80",  X"00",  X"2C",
  X"B0",  X"2C",  X"B8",  X"01",  X"E4",  X"00",  X"00",  X"08",
  X"00",  X"A0",  X"44",  X"44",  X"00",  X"00",  X"00",  X"44",
  X"00",  X"00",  X"44",  X"00",  X"40",  X"44",  X"00",  X"FF",
  X"0C",  X"05",  X"D0",  X"04",  X"AC",  X"00",  X"04",  X"1C",
  X"03",  X"A7",  X"00",  X"44",  X"00",  X"44",  X"00",  X"40",
  X"10",  X"40",  X"44",  X"00",  X"44",  X"00",  X"40",  X"08",
  X"40",  X"00",  X"08",  X"00",  X"A0",  X"44",  X"48",  X"44",
  X"00",  X"44",  X"00",  X"0C",  X"01",  X"48",  X"02",  X"02",
  X"02",  X"0C",  X"00",  X"08",  X"00",  X"A0",  X"44",  X"30",
  X"8C",  X"63",  X"00",  X"44",  X"04",  X"01",  X"76",  X"00",
  X"44",  X"01",  X"B7",  X"00",  X"00",  X"08",  X"00",  X"88",
  X"30",  X"84",  X"EB",  X"00",  X"2C",  X"70",  X"00",  X"F0",
  X"15",  X"FC",  X"00",  X"00",  X"08",  X"00",  X"00",  X"00",
  X"00",  X"2C",  X"00",  X"00",  X"D0",  X"08",  X"40",  X"FF",
  X"FF",  X"48",  X"3C",  X"FF",  X"44",  X"42",  X"18",  X"34",
  X"1A",  X"1B",  X"AD",  X"34",  X"34",  X"00",  X"08",  X"08",
  X"D0",  X"2D",  X"F0",  X"08",  X"40",  X"FF",  X"FF",  X"48",
  X"3C",  X"FF",  X"44",  X"34",  X"42",  X"19",  X"1A",  X"98",
  X"34",  X"34",  X"00",  X"08",  X"08",  X"A0",  X"31",  X"0C",
  X"9C",  X"2D",  X"28",  X"48",  X"00",  X"3D",  X"4C",  X"04",
  X"1F",  X"1E",  X"00",  X"00",  X"12",  X"02",  X"04",  X"22",
  X"42",  X"02",  X"02",  X"88",  X"04",  X"03",  X"01",  X"02",
  X"03",  X"88",  X"02",  X"19",  X"02",  X"02",  X"02",  X"01",
  X"04",  X"02",  X"00",  X"FE",  X"9C",  X"08",  X"00",  X"28",
  X"90",  X"00",  X"1A",  X"9C",  X"48",  X"00",  X"48",  X"04",
  X"88",  X"8C",  X"D9",  X"00",  X"8C",  X"03",  X"02",  X"02",
  X"02",  X"8C",  X"01",  X"02",  X"04",  X"00",  X"E3",  X"9C",
  X"08",  X"00",  X"C5",  X"48",  X"DD",  X"FF",  X"08",  X"00",
  X"08",  X"2D",  X"F0",  X"00",  X"18",  X"00",  X"00",  X"08",
  X"2D",  X"F0",  X"00",  X"03",  X"00",  X"00",  X"A0",  X"00",
  X"0B",  X"16",  X"04",  X"10",  X"F8",  X"1F",  X"19",  X"46",
  X"FF",  X"44",  X"00",  X"AF",  X"18",  X"F7",  X"41",  X"09",
  X"2F",  X"48",  X"10",  X"0C",  X"01",  X"0F",  X"03",  X"04",
  X"0C",  X"08",  X"FC",  X"03",  X"04",  X"01",  X"08",  X"04",
  X"0C",  X"18",  X"92",  X"08",  X"08",  X"00",  X"08",  X"04",
  X"FC",  X"10",  X"0F",  X"D2",  X"14",  X"31",  X"30",  X"10",
  X"54",  X"10",  X"FF",  X"04",  X"10",  X"FF",  X"00",  X"18",
  X"88",  X"15",  X"FF",  X"09",  X"08",  X"14",  X"08",  X"EC",
  X"31",  X"13",  X"EA",  X"1C",  X"08",  X"04",  X"FC",  X"10",
  X"0F",  X"22",  X"02",  X"69",  X"18",  X"08",  X"00",  X"03",
  X"00",  X"0F",  X"03",  X"04",  X"92",  X"06",  X"5B",  X"14",
  X"08",  X"03",  X"54",  X"13",  X"54",  X"0C",  X"6E",  X"03",
  X"2F",  X"48",  X"03",  X"0C",  X"12",  X"0B",  X"04",  X"10",
  X"01",  X"68",  X"0C",  X"0C",  X"12",  X"0A",  X"01",  X"04",
  X"FC",  X"10",  X"0F",  X"F6",  X"00",  X"FF",  X"01",  X"2F",
  X"50",  X"08",  X"12",  X"2A",  X"04",  X"04",  X"FC",  X"10",
  X"0F",  X"8A",  X"00",  X"0C",  X"59",  X"08",  X"FF",  X"62",
  X"03",  X"09",  X"04",  X"E9",  X"5B",  X"06",  X"38",  X"03",
  X"0D",  X"08",  X"0D",  X"08",  X"04",  X"E9",  X"04",  X"01",
  X"08",  X"0C",  X"04",  X"FC",  X"04",  X"FA",  X"08",  X"0C",
  X"0C",  X"08",  X"0C",  X"08",  X"04",  X"02",  X"01",  X"02",
  X"04",  X"7E",  X"08",  X"04",  X"4B",  X"FC",  X"03",  X"0C",
  X"0A",  X"0A",  X"0C",  X"12",  X"0B",  X"04",  X"58",  X"01",
  X"19",  X"0C",  X"0C",  X"12",  X"52",  X"01",  X"04",  X"FC",
  X"10",  X"0F",  X"F6",  X"00",  X"0C",  X"08",  X"10",  X"01",
  X"08",  X"0C",  X"0C",  X"08",  X"04",  X"01",  X"08",  X"10",
  X"0C",  X"08",  X"02",  X"04",  X"01",  X"08",  X"04",  X"0C",
  X"18",  X"DB",  X"08",  X"08",  X"00",  X"02",  X"04",  X"01",
  X"04",  X"18",  X"D2",  X"08",  X"08",  X"00",  X"38",  X"79",
  X"03",  X"03",  X"04",  X"08",  X"04",  X"0C",  X"08",  X"02",
  X"01",  X"0C",  X"02",  X"08",  X"0B",  X"B0",  X"04",  X"01",
  X"04",  X"FE",  X"04",  X"B4",  X"03",  X"31",  X"31",  X"08",
  X"10",  X"01",  X"01",  X"04",  X"04",  X"18",  X"08",  X"AD",
  X"08",  X"08",  X"00",  X"10",  X"BE",  X"01",  X"03",  X"A3",
  X"08",  X"03",  X"9C",  X"F8",  X"08",  X"01",  X"FB",  X"FF",
  X"04",  X"01",  X"01",  X"0B",  X"00",  X"0A",  X"08",  X"01",
  X"92",  X"01",  X"8C",  X"0B",  X"08",  X"0C",  X"12",  X"50",
  X"02",  X"EF",  X"04",  X"1C",  X"01",  X"12",  X"67",  X"1C",
  X"54",  X"FF",  X"6B",  X"30",  X"01",  X"02",  X"1C",  X"07",
  X"06",  X"04",  X"08",  X"02",  X"01",  X"00",  X"15",  X"18",
  X"FF",  X"15",  X"7E",  X"15",  X"FF",  X"60",  X"01",  X"12",
  X"15",  X"01",  X"1C",  X"01",  X"1C",  X"04",  X"13",  X"10",
  X"08",  X"0F",  X"3A",  X"F4",  X"F8",  X"02",  X"04",  X"01",
  X"04",  X"04",  X"05",  X"08",  X"0F",  X"42",  X"04",  X"31",
  X"14",  X"03",  X"02",  X"14",  X"31",  X"18",  X"03",  X"DD",
  X"18",  X"DC",  X"08",  X"95",  X"08",  X"DE",  X"17",  X"54",
  X"0F",  X"77",  X"EE",  X"03",  X"14",  X"1B",  X"03",  X"54",
  X"17",  X"54",  X"0C",  X"6E",  X"14",  X"03",  X"02",  X"01",
  X"04",  X"02",  X"04",  X"1D",  X"01",  X"F0",  X"DA",  X"7E",
  X"12",  X"7C",  X"D6",  X"03",  X"01",  X"B7",  X"04",  X"18",
  X"54",  X"0F",  X"77",  X"FD",  X"03",  X"FF",  X"9B",  X"54",
  X"08",  X"14",  X"01",  X"C4",  X"04",  X"9A",  X"54",  X"08",
  X"6C",  X"18",  X"31",  X"BC",  X"1C",  X"A5",  X"00",  X"F0",
  X"E8",  X"7E",  X"12",  X"7C",  X"E4",  X"03",  X"04",  X"04",
  X"68",  X"04",  X"6D",  X"04",  X"30",  X"58",  X"00",  X"12",
  X"00",  X"00",  X"30",  X"58",  X"00",  X"F6",  X"00",  X"00",
  X"A0",  X"32",  X"19",  X"93",  X"80",  X"FF",  X"04",  X"80",
  X"08",  X"08",  X"00",  X"FD",  X"00",  X"00",  X"08",  X"08",
  X"3C",  X"10",  X"10",  X"20",  X"10",  X"10",  X"10",  X"10",
  X"10",  X"10",  X"90",  X"3C",  X"10",  X"A4",  X"40",  X"10",
  X"4C",  X"5C",  X"5C",  X"5C",  X"5C",  X"5C",  X"5C",  X"5C",
  X"5C",  X"5C",  X"10",  X"10",  X"10",  X"10",  X"10",  X"10",
  X"10",  X"10",  X"10",  X"B4",  X"20",  X"6C",  X"10",  X"6C",
  X"10",  X"10",  X"10",  X"10",  X"5C",  X"10",  X"10",  X"D8",
  X"10",  X"10",  X"10",  X"AC",  X"10",  X"08",  X"10",  X"10",
  X"1C",  X"10",  X"10",  X"10",  X"10",  X"10",  X"10",  X"10",
  X"10",  X"10",  X"10",  X"B4",  X"24",  X"6C",  X"6C",  X"6C",
  X"9C",  X"24",  X"10",  X"10",  X"CC",  X"10",  X"FC",  X"DC",
  X"90",  X"BC",  X"10",  X"AC",  X"10",  X"0C",  X"10",  X"10",
  X"EC",  X"A0",  X"08",  X"00",  X"05",  X"18",  X"04",  X"08",
  X"00",  X"82",  X"19",  X"04",  X"08",  X"08",  X"08",  X"70",
  X"FA",  X"00",  X"00",  X"0C",  X"44",  X"00",  X"08",  X"E8",
  X"2D",  X"F0",  X"00",  X"07",  X"0C",  X"38",  X"00",  X"03",
  X"00",  X"0C",  X"08",  X"6E",  X"01",  X"10",  X"00",  X"6A",
  X"1A",  X"0A",  X"73",  X"0E",  X"40",  X"B4",  X"B0",  X"AC",
  X"F8",  X"FC",  X"EC",  X"F0",  X"2D",  X"2D",  X"A8",  X"98",
  X"00",  X"13",  X"00",  X"25",  X"1E",  X"00",  X"00",  X"1C",
  X"18",  X"1A",  X"01",  X"00",  X"25",  X"04",  X"00",  X"FC",
  X"01",  X"1A",  X"DE",  X"14",  X"04",  X"00",  X"08",  X"B0",
  X"B4",  X"01",  X"15",  X"B0",  X"07",  X"C1",  X"B4",  X"00",
  X"14",  X"15",  X"18",  X"00",  X"76",  X"01",  X"FF",  X"FF",
  X"00",  X"18",  X"00",  X"00",  X"2B",  X"20",  X"18",  X"01",
  X"E0",  X"58",  X"B9",  X"02",  X"00",  X"65",  X"01",  X"18",
  X"FF",  X"10",  X"08",  X"01",  X"18",  X"00",  X"02",  X"1A",
  X"84",  X"10",  X"02",  X"10",  X"17",  X"0C",  X"FF",  X"00",
  X"52",  X"02",  X"01",  X"04",  X"FF",  X"00",  X"B4",  X"B0",
  X"01",  X"01",  X"B0",  X"B4",  X"07",  X"57",  X"08",  X"0C",
  X"80",  X"5D",  X"10",  X"08",  X"1D",  X"00",  X"38",  X"10",
  X"24",  X"0C",  X"10",  X"10",  X"01",  X"06",  X"03",  X"F0",
  X"10",  X"19",  X"01",  X"04",  X"00",  X"08",  X"B0",  X"B4",
  X"01",  X"10",  X"B0",  X"07",  X"F3",  X"B4",  X"E4",  X"19",
  X"51",  X"AC",  X"00",  X"CB",  X"E4",  X"F0",  X"10",  X"EC",
  X"13",  X"01",  X"10",  X"02",  X"04",  X"0C",  X"00",  X"B4",
  X"01",  X"B4",  X"B0",  X"01",  X"B0",  X"07",  X"08",  X"08",
  X"19",  X"38",  X"AC",  X"00",  X"B2",  X"13",  X"00",  X"5B",
  X"65",  X"04",  X"00",  X"08",  X"B4",  X"1D",  X"B4",  X"B0",
  X"01",  X"07",  X"34",  X"B0",  X"04",  X"36",  X"B4",  X"10",
  X"01",  X"00",  X"30",  X"10",  X"1D",  X"04",  X"10",  X"06",
  X"AC",  X"F0",  X"10",  X"17",  X"04",  X"04",  X"00",  X"08",
  X"B0",  X"B4",  X"01",  X"10",  X"B0",  X"07",  X"F3",  X"B4",
  X"19",  X"08",  X"17",  X"00",  X"82",  X"F0",  X"10",  X"EE",
  X"13",  X"04",  X"04",  X"00",  X"B4",  X"01",  X"B0",  X"01",
  X"B4",  X"07",  X"09",  X"B0",  X"19",  X"F4",  X"AC",  X"00",
  X"6F",  X"00",  X"B4",  X"10",  X"03",  X"02",  X"03",  X"00",
  X"60",  X"1C",  X"B0",  X"00",  X"1E",  X"13",  X"44",  X"C5",
  X"16",  X"1A",  X"00",  X"08",  X"00",  X"01",  X"00",  X"00",
  X"32",  X"00",  X"10",  X"10",  X"2D",  X"00",  X"40",  X"2A",
  X"00",  X"02",  X"1D",  X"04",  X"00",  X"01",  X"FF",  X"00",
  X"02",  X"7F",  X"74",  X"00",  X"05",  X"DC",  X"FF",  X"3D",
  X"FF",  X"FF",  X"01",  X"33",  X"02",  X"26",  X"74",  X"07",
  X"FF",  X"30",  X"03",  X"00",  X"FB",  X"00",  X"DC",  X"01",
  X"33",  X"17",  X"30",  X"30",  X"30",  X"FF",  X"17",  X"2C",
  X"00",  X"1D",  X"04",  X"00",  X"DA",  X"01",  X"10",  X"10",
  X"0B",  X"00",  X"40",  X"08",  X"00",  X"02",  X"1D",  X"04",
  X"00",  X"CD",  X"00",  X"1D",  X"04",  X"00",  X"C8",  X"00",
  X"10",  X"10",  X"10",  X"40",  X"00",  X"04",  X"00",  X"52",
  X"1D",  X"01",  X"BD",  X"00",  X"06",  X"74",  X"01",  X"DF",
  X"30",  X"74",  X"00",  X"16",  X"03",  X"10",  X"10",  X"08",
  X"00",  X"FF",  X"00",  X"EC",  X"02",  X"10",  X"01",  X"10",
  X"84",  X"ED",  X"0C",  X"10",  X"02",  X"00",  X"E8",  X"10",
  X"24",  X"04",  X"10",  X"10",  X"01",  X"06",  X"03",  X"F0",
  X"10",  X"19",  X"01",  X"04",  X"00",  X"08",  X"B0",  X"B4",
  X"01",  X"10",  X"B0",  X"07",  X"F3",  X"B4",  X"E4",  X"19",
  X"51",  X"AC",  X"00",  X"CB",  X"E4",  X"F0",  X"10",  X"EC",
  X"13",  X"01",  X"10",  X"02",  X"04",  X"04",  X"00",  X"B4",
  X"01",  X"B4",  X"B0",  X"01",  X"B0",  X"07",  X"B8",  X"08",
  X"19",  X"38",  X"AC",  X"00",  X"B2",  X"FF",  X"00",  X"B3",
  X"13",  X"02",  X"BE",  X"0C",  X"F9",  X"30",  X"F8",  X"02",
  X"04",  X"F8",  X"00",  X"B4",  X"B0",  X"01",  X"02",  X"B0",
  X"B4",  X"07",  X"AD",  X"08",  X"19",  X"1C",  X"AC",  X"00",
  X"96",  X"0C",  X"80",  X"A8",  X"13",  X"10",  X"02",  X"00",
  X"A3",  X"10",  X"24",  X"0C",  X"10",  X"10",  X"01",  X"06",
  X"03",  X"F0",  X"10",  X"19",  X"01",  X"04",  X"00",  X"08",
  X"B0",  X"B4",  X"01",  X"10",  X"B0",  X"07",  X"F3",  X"B4",
  X"E4",  X"19",  X"F7",  X"AC",  X"00",  X"71",  X"E4",  X"F0",
  X"10",  X"EC",  X"13",  X"01",  X"10",  X"02",  X"04",  X"0C",
  X"00",  X"B4",  X"01",  X"B4",  X"B0",  X"01",  X"B0",  X"07",
  X"73",  X"08",  X"19",  X"DE",  X"AC",  X"00",  X"58",  X"13",
  X"6C",  X"08",  X"AC",  X"F4",  X"2D",  X"F8",  X"90",  X"00",
  X"48",  X"00",  X"F8",  X"F4",  X"01",  X"04",  X"2D",  X"78",
  X"B4",  X"00",  X"B0",  X"01",  X"01",  X"B0",  X"B4",  X"07",
  X"13",  X"08",  X"F4",  X"F4",  X"02",  X"06",  X"01",  X"01",
  X"95",  X"04",  X"01",  X"04",  X"E8",  X"00",  X"B0",  X"B4",
  X"01",  X"01",  X"B0",  X"B4",  X"07",  X"06",  X"08",  X"F4",
  X"FF",  X"00",  X"82",  X"10",  X"74",  X"0C",  X"10",  X"06",
  X"AC",  X"F0",  X"10",  X"6E",  X"04",  X"04",  X"00",  X"08",
  X"B0",  X"B4",  X"01",  X"10",  X"B0",  X"07",  X"F3",  X"B4",
  X"19",  X"90",  X"1D",  X"00",  X"0A",  X"13",  X"EC",  X"F0",
  X"19",  X"88",  X"AC",  X"00",  X"9F",  X"B0",  X"00",  X"06",
  X"0C",  X"44",  X"62",  X"16",  X"0C",  X"10",  X"10",  X"00",
  X"9E",  X"00",  X"40",  X"04",  X"00",  X"08",  X"00",  X"08",
  X"FF",  X"59",  X"19",  X"00",  X"1D",  X"0C",  X"0C",  X"03",
  X"1A",  X"0A",  X"93",  X"40",  X"0E",  X"00",  X"8E",  X"0E",
  X"00",  X"E6",  X"00",  X"FD",  X"24",  X"98",  X"18",  X"1C",
  X"84",  X"74",  X"00",  X"80",  X"82",  X"90",  X"80",  X"88",
  X"7C",  X"11",  X"FA",  X"8C",  X"11",  X"0D",  X"01",  X"11",
  X"CC",  X"BA",  X"10",  X"FC",  X"11",  X"44",  X"74",  X"1A",
  X"11",  X"4E",  X"1B",  X"00",  X"08",  X"80",  X"B8",  X"11",
  X"00",  X"02",  X"FF",  X"80",  X"40",  X"05",  X"00",  X"0C",
  X"40",  X"0C",  X"AE",  X"10",  X"08",  X"00",  X"01",  X"B6",
  X"01",  X"00",  X"F8",  X"2E",  X"F9",  X"02",  X"04",  X"F8",
  X"00",  X"B4",  X"B0",  X"01",  X"02",  X"B0",  X"B4",  X"07",
  X"BB",  X"08",  X"2D",  X"F8",  X"90",  X"00",  X"48",  X"00",
  X"72",  X"F4",  X"F4",  X"FF",  X"04",  X"01",  X"00",  X"B4",
  X"01",  X"B4",  X"B0",  X"01",  X"B0",  X"07",  X"9D",  X"08",
  X"F0",  X"04",  X"E0",  X"F0",  X"00",  X"B4",  X"B0",  X"01",
  X"03",  X"B4",  X"B0",  X"07",  X"D0",  X"08",  X"19",  X"F2",
  X"AC",  X"00",  X"6C",  X"13",  X"C9",  X"04",  X"19",  X"EA",
  X"AC",  X"00",  X"6A",  X"13",  X"3C",  X"00",  X"6D",  X"58",
  X"F9",  X"2D",  X"11",  X"00",  X"FE",  X"0C",  X"7B",  X"58",
  X"62",  X"0C",  X"00",  X"39",  X"F4",  X"02",  X"DD",  X"04",
  X"04",  X"F4",  X"00",  X"B0",  X"B4",  X"01",  X"03",  X"B0",
  X"B4",  X"07",  X"6F",  X"08",  X"F4",  X"F4",  X"01",  X"00",
  X"01",  X"10",  X"ED",  X"0C",  X"10",  X"06",  X"AC",  X"F0",
  X"10",  X"E7",  X"04",  X"04",  X"00",  X"08",  X"B0",  X"B4",
  X"01",  X"10",  X"B0",  X"07",  X"F3",  X"B4",  X"19",  X"AA",
  X"1D",  X"00",  X"24",  X"13",  X"EC",  X"F0",  X"73",  X"73",
  X"23",  X"01",  X"FF",  X"00",  X"9C",  X"10",  X"45",  X"0C",
  X"10",  X"06",  X"AC",  X"F0",  X"10",  X"3F",  X"04",  X"04",
  X"00",  X"08",  X"B0",  X"B4",  X"01",  X"10",  X"B0",  X"07",
  X"F3",  X"B4",  X"19",  X"86",  X"1D",  X"00",  X"00",  X"13",
  X"EC",  X"F0",  X"F3",  X"00",  X"02",  X"F1",  X"04",  X"1A",
  X"58",  X"0C",  X"19",  X"0E",  X"00",  X"00",  X"26",  X"04",
  X"1C",  X"00",  X"04",  X"D3",  X"18",  X"43",  X"23",  X"10",
  X"22",  X"D8",  X"00",  X"01",  X"04",  X"18",  X"18",  X"1D",
  X"FF",  X"1F",  X"08",  X"01",  X"00",  X"D1",  X"10",  X"10",
  X"C0",  X"00",  X"40",  X"BD",  X"00",  X"04",  X"8C",  X"00",
  X"00",  X"01",  X"B4",  X"18",  X"00",  X"B1",  X"18",  X"FF",
  X"00",  X"AD",  X"18",  X"00",  X"80",  X"A9",  X"18",  X"D0",
  X"00",  X"00",  X"03",  X"01",  X"02",  X"1C",  X"D0",  X"09",
  X"F9",  X"01",  X"9F",  X"E0",  X"00",  X"1D",  X"2D",  X"04",
  X"58",  X"00",  X"02",  X"EC",  X"02",  X"61",  X"78",  X"00",
  X"10",  X"8D",  X"18",  X"00",  X"18",  X"18",  X"6C",  X"04",
  X"01",  X"85",  X"10",  X"2D",  X"58",  X"10",  X"4E",  X"EC",
  X"40",  X"4C",  X"00",  X"02",  X"04",  X"1D",  X"00",  X"00",
  X"46",  X"02",  X"01",  X"44",  X"FF",  X"02",  X"40",  X"01",
  X"00",  X"2A",  X"48",  X"01",  X"D0",  X"00",  X"09",  X"69",
  X"00",  X"00",  X"03",  X"01",  X"0D",  X"01",  X"D0",  X"09",
  X"F9",  X"01",  X"00",  X"5D",  X"FF",  X"5C",  X"E0",  X"00",
  X"40",  X"55",  X"18",  X"FF",  X"00",  X"00",  X"73",  X"04",
  X"53",  X"C7",  X"10",  X"C6",  X"F0",  X"00",  X"AB",  X"17",
  X"00",  X"67",  X"16",  X"00",  X"07",  X"10",  X"17",  X"16",
  X"3B",  X"1D",  X"10",  X"16",  X"08",  X"5C",  X"00",  X"2D",
  X"38",  X"10",  X"B6",  X"EC",  X"00",  X"B8",  X"04",  X"FF",
  X"00",  X"7C",  X"00",  X"FF",  X"00",  X"29",  X"18",  X"00",
  X"08",  X"25",  X"18",  X"FF",  X"9D",  X"47",  X"08",  X"67",
  X"07",  X"00",  X"08",  X"8D",  X"1B",  X"C8",  X"76",  X"08",
  X"C8",  X"F8",  X"10",  X"08",  X"82",  X"F8",  X"00",  X"90",
  X"2D",  X"F8",  X"90",  X"00",  X"C8",  X"00",  X"FD",  X"2D",
  X"03",  X"2D",  X"10",  X"03",  X"08",  X"50",  X"23",  X"00",
  X"04",  X"D1",  X"00",  X"EC",  X"0F",  X"01",  X"FF",  X"04",
  X"00",  X"FB",  X"00",  X"DC",  X"0F",  X"17",  X"09",  X"10",
  X"74",  X"02",  X"1D",  X"0A",  X"DF",  X"FF",  X"30",  X"0A",
  X"1D",  X"2E",  X"00",  X"09",  X"F6",  X"08",  X"17",  X"30",
  X"DC",  X"FF",  X"FF",  X"F8",  X"17",  X"4D",  X"00",  X"01",
  X"04",  X"00",  X"08",  X"B0",  X"B4",  X"01",  X"01",  X"B0",
  X"07",  X"67",  X"B4",  X"19",  X"65",  X"AC",  X"00",  X"DF",
  X"13",  X"60",  X"F0",  X"19",  X"5D",  X"AC",  X"00",  X"D7",
  X"13",  X"42",  X"2D",  X"04",  X"0C",  X"00",  X"B4",  X"15",
  X"B0",  X"01",  X"B4",  X"B0",  X"07",  X"4B",  X"08",  X"E5",
  X"19",  X"D8",  X"00",  X"08",  X"9B",  X"16",  X"00",  X"44",
  X"16",  X"18",  X"AD",  X"17",  X"FF",  X"28",  X"08",  X"D8",
  X"04",  X"2D",  X"1D",  X"FF",  X"1D",  X"01",  X"69",  X"00",
  X"04",  X"0C",  X"00",  X"B4",  X"15",  X"08",  X"01",  X"B4",
  X"C0",  X"EB",  X"08",  X"C0",  X"F8",  X"08",  X"76",  X"10",
  X"F0",  X"00",  X"D0",  X"74",  X"08",  X"00",  X"F4",  X"00",
  X"00",  X"10",  X"15",  X"10",  X"1D",  X"16",  X"03",  X"01",
  X"01",  X"F0",  X"16",  X"00",  X"C4",  X"44",  X"18",  X"78",
  X"D0",  X"FF",  X"F4",  X"0C",  X"10",  X"1D",  X"BA",  X"01",
  X"F0",  X"04",  X"15",  X"1B",  X"10",  X"00",  X"92",  X"00",
  X"10",  X"80",  X"08",  X"00",  X"08",  X"B4",  X"01",  X"B4",
  X"B0",  X"01",  X"07",  X"A6",  X"B0",  X"01",  X"F4",  X"04",
  X"2D",  X"80",  X"B4",  X"00",  X"B0",  X"01",  X"01",  X"B0",
  X"B4",  X"07",  X"8F",  X"08",  X"F4",  X"F4",  X"01",  X"04",
  X"15",  X"00",  X"B4",  X"01",  X"B0",  X"DB",  X"01",  X"04",
  X"0C",  X"00",  X"B4",  X"15",  X"B0",  X"01",  X"B4",  X"B0",
  X"07",  X"08",  X"08",  X"19",  X"C5",  X"AC",  X"00",  X"3F",
  X"13",  X"01",  X"9B",  X"04",  X"01",  X"04",  X"2D",  X"80",
  X"B4",  X"00",  X"B0",  X"01",  X"BD",  X"01",  X"00",  X"FB",
  X"01",  X"FA",  X"08",  X"19",  X"AD",  X"AC",  X"00",  X"27",
  X"13",  X"EA",  X"F4",  X"04",  X"2D",  X"FF",  X"10",  X"03",
  X"50",  X"08",  X"2E",  X"00",  X"01",  X"04",  X"2D",  X"78",
  X"B4",  X"00",  X"B0",  X"01",  X"01",  X"B0",  X"B4",  X"07",
  X"51",  X"08",  X"F4",  X"00",  X"30",  X"F4",  X"01",  X"04",
  X"E8",  X"00",  X"B0",  X"B4",  X"01",  X"01",  X"B0",  X"B4",
  X"07",  X"64",  X"08",  X"F4",  X"15",  X"00",  X"F5",  X"10",
  X"E1",  X"0C",  X"10",  X"06",  X"AC",  X"F0",  X"10",  X"DB",
  X"04",  X"04",  X"00",  X"08",  X"B0",  X"B4",  X"01",  X"10",
  X"B0",  X"07",  X"F3",  X"B4",  X"19",  X"64",  X"10",  X"00",
  X"DE",  X"13",  X"EC",  X"F0",  X"00",  X"38",  X"04",  X"D0",
  X"01",  X"19",  X"57",  X"AC",  X"00",  X"D1",  X"13",  X"8E",
  X"F4",  X"19",  X"4F",  X"AC",  X"00",  X"C9",  X"13",  X"6E",
  X"F4",  X"19",  X"47",  X"AC",  X"00",  X"C1",  X"13",  X"57",
  X"01",  X"19",  X"3F",  X"AC",  X"00",  X"B9",  X"13",  X"AC",
  X"F4",  X"08",  X"A4",  X"00",  X"08",  X"08",  X"1F",  X"01",
  X"B9",  X"10",  X"B4",  X"00",  X"05",  X"19",  X"B0",  X"AE",
  X"0C",  X"28",  X"AC",  X"00",  X"A9",  X"0C",  X"B0",  X"A6",
  X"0C",  X"69",  X"06",  X"00",  X"10",  X"81",  X"18",  X"FC",
  X"F8",  X"00",  X"A7",  X"03",  X"00",  X"66",  X"16",  X"07",
  X"03",  X"45",  X"00",  X"65",  X"FE",  X"02",  X"F8",  X"B8",
  X"0C",  X"B8",  X"00",  X"1D",  X"28",  X"EC",  X"44",  X"5C",
  X"10",  X"E8",  X"14",  X"60",  X"1D",  X"B8",  X"F4",  X"47",
  X"C2",  X"08",  X"67",  X"C0",  X"01",  X"2D",  X"66",  X"1D",
  X"0E",  X"90",  X"00",  X"10",  X"48",  X"00",  X"B9",  X"E8",
  X"E8",  X"67",  X"17",  X"01",  X"FF",  X"47",  X"05",  X"F4",
  X"00",  X"9C",  X"65",  X"F4",  X"FD",  X"06",  X"00",  X"1D",
  X"9A",  X"F4",  X"00",  X"45",  X"04",  X"45",  X"65",  X"65",
  X"FF",  X"E0",  X"00",  X"08",  X"F4",  X"2B",  X"E1",  X"09",
  X"BD",  X"A8",  X"30",  X"30",  X"E2",  X"E3",  X"E4",  X"F4",
  X"01",  X"E0",  X"01",  X"F4",  X"F0",  X"11",  X"02",  X"01",
  X"0C",  X"FF",  X"19",  X"1D",  X"2D",  X"08",  X"FF",  X"00",
  X"1D",  X"1F",  X"01",  X"01",  X"3C",  X"10",  X"01",  X"F2",
  X"0C",  X"F0",  X"01",  X"19",  X"A5",  X"AC",  X"00",  X"1F",
  X"13",  X"F7",  X"F4",  X"08",  X"1F",  X"00",  X"01",  X"22",
  X"10",  X"04",  X"0C",  X"00",  X"B4",  X"15",  X"B0",  X"01",
  X"B4",  X"B0",  X"07",  X"08",  X"08",  X"19",  X"8B",  X"AC",
  X"00",  X"05",  X"13",  X"F4",  X"04",  X"00",  X"08",  X"B4",
  X"B0",  X"01",  X"03",  X"B0",  X"07",  X"57",  X"B4",  X"88",
  X"19",  X"06",  X"2D",  X"10",  X"06",  X"88",  X"08",  X"E7",
  X"00",  X"2D",  X"10",  X"03",  X"08",  X"70",  X"F3",  X"00",
  X"44",  X"3D",  X"01",  X"00",  X"51",  X"08",  X"00",  X"B8",
  X"D0",  X"44",  X"16",  X"D0",  X"F0",  X"ED",  X"1D",  X"08",
  X"B8",  X"1D",  X"1D",  X"16",  X"1F",  X"08",  X"01",  X"DA",
  X"10",  X"00",  X"DD",  X"58",  X"ED",  X"FF",  X"08",  X"00",
  X"10",  X"15",  X"1B",  X"4A",  X"10",  X"58",  X"66",  X"8B",
  X"F4",  X"F4",  X"1D",  X"63",  X"00",  X"01",  X"82",  X"67",
  X"80",  X"01",  X"01",  X"43",  X"2D",  X"4C",  X"E8",  X"04",
  X"04",  X"8D",  X"30",  X"00",  X"01",  X"01",  X"FD",  X"E8",
  X"42",  X"67",  X"44",  X"00",  X"F0",  X"00",  X"B4",  X"D0",
  X"FF",  X"0C",  X"08",  X"22",  X"F0",  X"19",  X"1B",  X"AC",
  X"00",  X"95",  X"13",  X"99",  X"F4",  X"0C",  X"40",  X"02",
  X"95",  X"0C",  X"01",  X"03",  X"02",  X"01",  X"E4",  X"1D",
  X"0A",  X"64",  X"FF",  X"30",  X"0A",  X"1D",  X"B3",  X"00",
  X"E4",  X"09",  X"F4",  X"08",  X"30",  X"FF",  X"16",  X"FF",
  X"02",  X"06",  X"E2",  X"35",  X"F4",  X"00",  X"01",  X"00",
  X"03",  X"FC",  X"01",  X"2D",  X"F4",  X"F4",  X"1A",  X"15",
  X"29",  X"AA",  X"2D",  X"10",  X"E1",  X"0C",  X"00",  X"30",
  X"0E",  X"2D",  X"F4",  X"1D",  X"EE",  X"90",  X"02",  X"03",
  X"1D",  X"01",  X"F4",  X"01",  X"1C",  X"67",  X"2D",  X"10",
  X"90",  X"00",  X"48",  X"00",  X"0B",  X"03",  X"01",  X"1D",
  X"F4",  X"D9",  X"1D",  X"2D",  X"1D",  X"FA",  X"E1",  X"F4",
  X"D2",  X"1D",  X"00",  X"00",  X"70",  X"04",  X"00",  X"18",
  X"1E",  X"FF",  X"00",  X"0B",  X"00",  X"06",  X"01",  X"01",
  X"F9",  X"0C",  X"01",  X"66",  X"F4",  X"16",  X"06",  X"02",
  X"01",  X"EF",  X"01",  X"02",  X"EC",  X"66",  X"BB",  X"04",
  X"0C",  X"40",  X"1F",  X"0C",  X"2D",  X"08",  X"F0",  X"09",
  X"0A",  X"02",  X"01",  X"00",  X"A3",  X"00",  X"00",  X"90",
  X"00",  X"0F",  X"18",  X"19",  X"1A",  X"18",  X"77",  X"1B",
  X"FF",  X"05",  X"08",  X"00",  X"8A",  X"00",  X"08",  X"00",
  X"18",  X"F0",  X"00",  X"6A",  X"1B",  X"F4",  X"FF",  X"2D",
  X"08",  X"F0",  X"09",  X"0A",  X"02",  X"01",  X"00",  X"E0",
  X"00",  X"00",  X"90",  X"00",  X"49",  X"18",  X"00",  X"3D",
  X"00",  X"00",  X"F0",  X"00",  X"04",  X"10",  X"11",  X"1C",
  X"CF",  X"19",  X"FF",  X"29",  X"00",  X"08",  X"18",  X"2A",
  X"04",  X"1B",  X"27",  X"04",  X"00",  X"0F",  X"08",  X"00",
  X"09",  X"00",  X"01",  X"01",  X"01",  X"01",  X"FD",  X"01",
  X"08",  X"00",  X"04",  X"00",  X"00",  X"00",  X"19",  X"1B",
  X"12",  X"04",  X"00",  X"00",  X"04",  X"10",  X"11",  X"A8",
  X"1C",  X"FF",  X"DC",  X"08",  X"8A",  X"00",  X"00",  X"08",
  X"FF",  X"00",  X"08",  X"00",  X"00",  X"08",  X"00",  X"00",
  X"02",  X"00",  X"00",  X"08",  X"FF",  X"00",  X"BB",  X"FF",
  X"2D",  X"08",  X"09",  X"F0",  X"0A",  X"0B",  X"03",  X"02",
  X"01",  X"00",  X"A8",  X"00",  X"00",  X"A0",  X"30",  X"7F",
  X"48",  X"01",  X"27",  X"48",  X"2D",  X"3F",  X"B8",  X"00",
  X"12",  X"00",  X"22",  X"7F",  X"1B",  X"00",  X"80",  X"7F",
  X"1E",  X"3F",  X"C0",  X"80",  X"06",  X"C0",  X"01",  X"00",
  X"08",  X"02",  X"48",  X"2D",  X"28",  X"C0",  X"00",  X"58",
  X"00",  X"0B",  X"08",  X"FF",  X"41",  X"20",  X"00",  X"08",
  X"01",  X"00",  X"FD",  X"00",  X"08",  X"00",  X"00",  X"3D",
  X"FF",  X"01",  X"74",  X"C0",  X"BF",  X"02",  X"FF",  X"01",
  X"12",  X"3F",  X"12",  X"80",  X"07",  X"0C",  X"F0",  X"3F",
  X"C0",  X"80",  X"06",  X"80",  X"03",  X"00",  X"01",  X"02",
  X"08",  X"04",  X"00",  X"FF",  X"02",  X"FF",  X"01",  X"6E",
  X"3F",  X"18",  X"80",  X"03",  X"12",  X"F8",  X"3F",  X"0C",
  X"80",  X"3F",  X"C0",  X"80",  X"06",  X"80",  X"04",  X"00",
  X"01",  X"02",  X"03",  X"08",  X"05",  X"FF",  X"0F",  X"50",
  X"7F",  X"80",  X"FF",  X"7C",  X"07",  X"1A",  X"C0",  X"FF",
  X"3E",  X"33",  X"FF",  X"01",  X"00",  X"08",  X"02",  X"48",
  X"2D",  X"CB",  X"C8",  X"00",  X"0E",  X"00",  X"AE",  X"08",
  X"FF",  X"A6",  X"00",  X"5F",  X"FF",  X"5D",  X"6C",  X"5F",
  X"08",  X"FF",  X"48",  X"2D",  X"B8",  X"D0",  X"00",  X"9B",
  X"00",  X"13",  X"01",  X"08",  X"FF",  X"41",  X"1A",  X"00",
  X"00",  X"0A",  X"1B",  X"00",  X"00",  X"28",  X"04",  X"01",
  X"42",  X"02",  X"03",  X"00",  X"08",  X"00",  X"CA",  X"01",
  X"FF",  X"DF",  X"3F",  X"0C",  X"80",  X"0F",  X"C0",  X"E0",
  X"06",  X"80",  X"02",  X"00",  X"01",  X"08",  X"03",  X"FF",
  X"1E",  X"B1",  X"80",  X"08",  X"FF",  X"3F",  X"1E",  X"80",
  X"01",  X"18",  X"FC",  X"3F",  X"12",  X"80",  X"3F",  X"0C",
  X"80",  X"3F",  X"C0",  X"80",  X"06",  X"80",  X"05",  X"00",
  X"01",  X"02",  X"03",  X"04",  X"08",  X"06",  X"DF",  X"FF",
  X"5D",  X"CB",  X"FF",  X"DF",  X"FF",  X"5D",  X"12",  X"00",
  X"00",  X"00",  X"0C",  X"02",  X"01",  X"00",  X"1B",  X"00",
  X"24",  X"05",  X"01",  X"42",  X"02",  X"03",  X"01",  X"00",
  X"08",  X"00",  X"FF",  X"5D",  X"B0",  X"FF",  X"01",  X"00",
  X"08",  X"02",  X"A0",  X"2D",  X"F0",  X"00",  X"06",  X"18",
  X"38",  X"00",  X"20",  X"00",  X"0C",  X"10",  X"10",  X"08",
  X"22",  X"01",  X"10",  X"00",  X"1A",  X"00",  X"0C",  X"01",
  X"0C",  X"02",  X"06",  X"00",  X"08",  X"00",  X"08",  X"00",
  X"14",  X"08",  X"08",  X"00",  X"14",  X"01",  X"08",  X"18",
  X"08",  X"00",  X"21",  X"00",  X"E1",  X"0C",  X"1A",  X"10",
  X"E7",  X"0C",  X"10",  X"EB",  X"FF",  X"04",  X"06",  X"30",
  X"08",  X"10",  X"D9",  X"0C",  X"00",  X"0B",  X"DB",  X"40",
  X"02",  X"07",  X"30",  X"B9",  X"F0",  X"0C",  X"30",  X"DB",
  X"10",  X"04",  X"0C",  X"08",  X"00",  X"C6",  X"0C",  X"A0",
  X"10",  X"10",  X"18",  X"01",  X"7F",  X"00",  X"03",  X"02",
  X"1D",  X"1D",  X"04",  X"04",  X"01",  X"1A",  X"69",  X"FF",
  X"04",  X"00",  X"14",  X"3B",  X"14",  X"3F",  X"11",  X"FF",
  X"1C",  X"00",  X"00",  X"00",  X"15",  X"20",  X"18",  X"10",
  X"08",  X"1C",  X"18",  X"00",  X"10",  X"15",  X"01",  X"15",
  X"10",  X"02",  X"08",  X"10",  X"15",  X"04",  X"01",  X"02",
  X"04",  X"00",  X"14",  X"04",  X"10",  X"E6",  X"10",  X"00",
  X"17",  X"19",  X"04",  X"02",  X"02",  X"01",  X"11",  X"10",
  X"02",  X"00",  X"08",  X"FC",  X"0B",  X"10",  X"00",  X"00",
  X"05",  X"FC",  X"01",  X"FB",  X"FF",  X"10",  X"19",  X"6C",
  X"10",  X"00",  X"31",  X"3F",  X"01",  X"FF",  X"1C",  X"00",
  X"00",  X"00",  X"10",  X"10",  X"0B",  X"02",  X"0B",  X"04",
  X"0C",  X"10",  X"04",  X"02",  X"04",  X"00",  X"11",  X"04",
  X"F0",  X"10",  X"04",  X"02",  X"02",  X"04",  X"00",  X"14",
  X"01",  X"12",  X"10",  X"02",  X"00",  X"0A",  X"FC",  X"10",
  X"08",  X"00",  X"00",  X"00",  X"07",  X"10",  X"FC",  X"01",
  X"FA",  X"FF",  X"10",  X"08",  X"00",  X"60",  X"40",  X"C8",
  X"CC",  X"00",  X"5C",  X"60",  X"10",  X"C8",  X"44",  X"04",
  X"01",  X"D4",  X"44",  X"02",  X"08",  X"D0",  X"01",  X"BF",
  X"18",  X"D0",  X"40",  X"D4",  X"C4",  X"C4",  X"00",  X"3E",
  X"01",  X"00",  X"00",  X"01",  X"01",  X"23",  X"2D",  X"28",
  X"90",  X"29",  X"4C",  X"00",  X"37",  X"01",  X"00",  X"2D",
  X"00",  X"15",  X"78",  X"2D",  X"79",  X"00",  X"08",  X"FF",
  X"01",  X"00",  X"EC",  X"18",  X"9A",  X"14",  X"00",  X"00",
  X"15",  X"EC",  X"01",  X"03",  X"00",  X"00",  X"08",  X"00",
  X"C4",  X"09",  X"0F",  X"00",  X"C4",  X"00",  X"FA",  X"00",
  X"2D",  X"70",  X"00",  X"08",  X"00",  X"03",  X"00",  X"03",
  X"03",  X"08",  X"00",  X"08",  X"00",  X"00",  X"00",  X"01",
  X"C4",  X"C1",  X"C4",  X"C8",  X"D4",  X"D0",  X"DC",  X"D8",
  X"18",  X"F8",  X"C8",  X"0C",  X"0D",  X"BB",  X"FC",  X"14",
  X"08",  X"FF",  X"D4",  X"D0",  X"DC",  X"D9",  X"D8",  X"C4",
  X"FC",  X"F8",  X"03",  X"32",  X"04",  X"20",  X"C4",  X"07",
  X"02",  X"12",  X"04",  X"03",  X"02",  X"03",  X"C4",  X"00",
  X"C4",  X"69",  X"0E",  X"C8",  X"CD",  X"C8",  X"0D",  X"00",
  X"0C",  X"02",  X"01",  X"E8",  X"C8",  X"C4",  X"2D",  X"F0",
  X"2D",  X"C8",  X"CE",  X"F8",  X"4C",  X"C4",  X"0D",  X"2D",
  X"00",  X"4C",  X"2D",  X"08",  X"4C",  X"4C",  X"90",  X"CE",
  X"4C",  X"C4",  X"00",  X"07",  X"C4",  X"0E",  X"4C",  X"00",
  X"02",  X"FF",  X"01",  X"16",  X"0B",  X"F4",  X"03",  X"2D",
  X"80",  X"02",  X"CC",  X"00",  X"03",  X"F4",  X"FF",  X"FF",
  X"00",  X"04",  X"00",  X"04",  X"01",  X"01",  X"00",  X"00",
  X"D9",  X"13",  X"E4",  X"F0",  X"13",  X"09",  X"8C",  X"FF",
  X"05",  X"04",  X"01",  X"FC",  X"00",  X"03",  X"0A",  X"00",
  X"D3",  X"02",  X"04",  X"1B",  X"05",  X"D0",  X"FF",  X"01",
  X"1C",  X"01",  X"00",  X"48",  X"E0",  X"44",  X"17",  X"01",
  X"D5",  X"04",  X"02",  X"01",  X"14",  X"04",  X"FC",  X"01",
  X"0F",  X"44",  X"00",  X"D4",  X"12",  X"D0",  X"DC",  X"D8",
  X"06",  X"18",  X"40",  X"08",  X"FF",  X"D4",  X"D0",  X"DC",
  X"70",  X"D8",  X"0E",  X"CC",  X"F8",  X"00",  X"C9",  X"2D",
  X"03",  X"00",  X"80",  X"6D",  X"01",  X"CC",  X"01",  X"01",
  X"4A",  X"C4",  X"0A",  X"4C",  X"CE",  X"C4",  X"30",  X"21",
  X"00",  X"2D",  X"18",  X"4A",  X"90",  X"4A",  X"00",  X"27",
  X"01",  X"18",  X"09",  X"90",  X"00",  X"4A",  X"00",  X"4A",
  X"00",  X"12",  X"EC",  X"CC",  X"01",  X"01",  X"4A",  X"C4",
  X"0A",  X"4C",  X"CE",  X"C4",  X"30",  X"00",  X"EE",  X"01",
  X"48",  X"C8",  X"00",  X"26",  X"FF",  X"48",  X"00",  X"FC",
  X"EC",  X"C4",  X"C4",  X"01",  X"1D",  X"FF",  X"F5",  X"EC",
  X"2D",  X"01",  X"08",  X"D8",  X"05",  X"2D",  X"C8",  X"00",
  X"01",  X"E8",  X"C8",  X"0C",  X"0D",  X"00",  X"0D",  X"01",
  X"3C",  X"FC",  X"E0",  X"00",  X"00",  X"01",  X"FF",  X"00",
  X"44",  X"00",  X"D4",  X"D0",  X"DC",  X"D8",  X"98",  X"18",
  X"40",  X"08",  X"FF",  X"D4",  X"D0",  X"DC",  X"94",  X"D8",
  X"00",  X"2F",  X"0F",  X"03",  X"2D",  X"2A",  X"80",  X"2B",
  X"01",  X"04",  X"10",  X"2A",  X"02",  X"00",  X"0E",  X"C8",
  X"2D",  X"48",  X"01",  X"05",  X"01",  X"00",  X"4E",  X"01",
  X"00",  X"F9",  X"08",  X"C8",  X"F4",  X"00",  X"20",  X"C4",
  X"2D",  X"10",  X"CC",  X"00",  X"19",  X"00",  X"00",  X"16",
  X"E0",  X"00",  X"D4",  X"01",  X"C4",  X"2D",  X"18",  X"4C",
  X"2D",  X"C4",  X"0C",  X"4E",  X"20",  X"4C",  X"C8",  X"00",
  X"C8",  X"0C",  X"FF",  X"63",  X"EC",  X"C4",  X"2D",  X"00",
  X"C4",  X"0C",  X"48",  X"20",  X"4C",  X"C8",  X"00",  X"C8",
  X"54",  X"0C",  X"C8",  X"2D",  X"28",  X"CC",  X"C8",  X"CC",
  X"00",  X"C3",  X"EC",  X"AC",  X"CC",  X"00",  X"A8",  X"00",
  X"EC",  X"00",  X"1C",  X"EC",  X"15",  X"0E",  X"00",  X"00",
  X"1D",  X"01",  X"F0",  X"E8",  X"EC",  X"00",  X"0D",  X"E8",
  X"00",  X"0A",  X"0C",  X"03",  X"1A",  X"0C",  X"E8",  X"01",
  X"E8",  X"01",  X"01",  X"F0",  X"00",  X"1B",  X"00",  X"4D",
  X"00",  X"13",  X"EC",  X"D4",  X"D0",  X"11",  X"0B",  X"18",
  X"EC",  X"14",  X"18",  X"3B",  X"EC",  X"14",  X"08",  X"DF",
  X"18",  X"D0",  X"D4",  X"12",  X"F0",  X"11",  X"52",  X"14",
  X"D4",  X"D0",  X"18",  X"B3",  X"01",  X"E4",  X"08",  X"00",
  X"D4",  X"09",  X"D0",  X"08",  X"03",  X"EC",  X"18",  X"D0",
  X"D4",  X"08",  X"01",  X"3A",  X"C4",  X"F0",  X"E4",  X"00",
  X"E9",  X"01",  X"1A",  X"1F",  X"70",  X"1C",  X"E8",  X"02",
  X"E8",  X"02",  X"02",  X"00",  X"0A",  X"14",  X"D4",  X"D0",
  X"19",  X"B8",  X"18",  X"D0",  X"D4",  X"08",  X"00",  X"0A",
  X"11",  X"D4",  X"D0",  X"1A",  X"AD",  X"18",  X"D0",  X"D4",
  X"08",  X"F4",  X"00",  X"D3",  X"D4",  X"00",  X"00",  X"02",
  X"00",  X"15",  X"77",  X"01",  X"E8",  X"00",  X"0A",  X"EC",
  X"D4",  X"D0",  X"0C",  X"96",  X"18",  X"D0",  X"EC",  X"D4",
  X"F0",  X"00",  X"34",  X"EC",  X"C4",  X"EC",  X"15",  X"01",
  X"C4",  X"01",  X"11",  X"24",  X"14",  X"30",  X"1C",  X"F4",
  X"DB",  X"14",  X"11",  X"F0",  X"17",  X"0F",  X"18",  X"0C",
  X"00",  X"08",  X"07",  X"01",  X"DC",  X"01",  X"68",  X"18",
  X"DC",  X"00",  X"08",  X"F0",  X"00",  X"06",  X"00",  X"00",
  X"33",  X"F4",  X"00",  X"E5",  X"00",  X"08",  X"00",  X"00",
  X"05",  X"00",  X"00",  X"DD",  X"00",  X"1A",  X"F4",  X"16",
  X"00",  X"3C",  X"01",  X"14",  X"18",  X"0A",  X"31",  X"00",
  X"17",  X"06",  X"08",  X"1C",  X"0A",  X"00",  X"29",  X"18",
  X"17",  X"08",  X"0A",  X"18",  X"00",  X"22",  X"01",  X"BB",
  X"08",  X"13",  X"F0",  X"2A",  X"E4",  X"2D",  X"68",  X"CC",
  X"0F",  X"D4",  X"03",  X"52",  X"FF",  X"00",  X"01",  X"E0",
  X"FF",  X"AF",  X"00",  X"18",  X"0A",  X"00",  X"09",  X"01",
  X"08",  X"11",  X"C5",  X"14",  X"30",  X"F4",  X"16",  X"00",
  X"14",  X"F2",  X"01",  X"EC",  X"00",  X"14",  X"01",  X"1A",
  X"18",  X"11",  X"71",  X"08",  X"00",  X"04",  X"FF",  X"A5",
  X"FF",  X"39",  X"FF",  X"B0",  X"FF",  X"15",  X"FA",  X"01",
  X"31",  X"00",  X"01",  X"11",  X"FA",  X"18",  X"00",  X"67",
  X"17",  X"06",  X"00",  X"04",  X"1C",  X"F1",  X"18",  X"17",
  X"EC",  X"ED",  X"18",  X"51",  X"18",  X"6B",  X"F0",  X"FF",
  X"01",  X"09",  X"01",  X"E4",  X"0D",  X"01",  X"01",  X"F0",
  X"E4",  X"00",  X"16",  X"E8",  X"00",  X"04",  X"00",  X"E8",
  X"16",  X"D4",  X"D0",  X"01",  X"01",  X"18",  X"B0",  X"01",
  X"D0",  X"EC",  X"CB",  X"D4",  X"EC",  X"16",  X"00",  X"AD",
  X"48",  X"FF",  X"03",  X"2D",  X"80",  X"01",  X"2D",  X"30",
  X"CC",  X"48",  X"C4",  X"0C",  X"CC",  X"C4",  X"30",  X"00",
  X"C8",  X"C8",  X"C8",  X"CC",  X"00",  X"16",  X"01",  X"2D",
  X"10",  X"CC",  X"CE",  X"00",  X"D3",  X"01",  X"40",  X"2D",
  X"10",  X"18",  X"0A",  X"01",  X"00",  X"CC",  X"C8",  X"00",
  X"28",  X"EC",  X"35",  X"2A",  X"50",  X"4C",  X"C4",  X"0E",
  X"CE",  X"50",  X"01",  X"C8",  X"02",  X"C4",  X"30",  X"00",
  X"00",  X"EB",  X"01",  X"F1",  X"18",  X"C4",  X"00",  X"C7",
  X"F0",  X"C4",  X"00",  X"C4",  X"02",  X"C1",  X"F0",  X"00",
  X"02",  X"BD",  X"F0",  X"01",  X"01",  X"01",  X"B8",  X"F0",
  X"FF",  X"39",  X"FF",  X"D5",  X"FF",  X"15",  X"FA",  X"01",
  X"30",  X"01",  X"00",  X"31",  X"CD",  X"15",  X"2A",  X"93",
  X"2B",  X"01",  X"DC",  X"C8",  X"14",  X"DC",  X"F6",  X"08",
  X"00",  X"95",  X"CC",  X"00",  X"4C",  X"2D",  X"28",  X"4A",
  X"C8",  X"00",  X"47",  X"EC",  X"00",  X"EC",  X"31",  X"01",
  X"00",  X"01",  X"51",  X"00",  X"20",  X"01",  X"04",  X"33",
  X"E8",  X"FC",  X"01",  X"01",  X"01",  X"8E",  X"E8",  X"1C",
  X"18",  X"0A",  X"00",  X"24",  X"01",  X"08",  X"BC",  X"08",
  X"2A",  X"2B",  X"13",  X"E9",  X"02",  X"0F",  X"2D",  X"03",
  X"80",  X"02",  X"04",  X"48",  X"00",  X"DF",  X"02",  X"2D",
  X"48",  X"01",  X"05",  X"01",  X"00",  X"4C",  X"01",  X"00",
  X"F9",  X"08",  X"D3",  X"F4",  X"C4",  X"0C",  X"CC",  X"01",
  X"01",  X"C4",  X"30",  X"2D",  X"80",  X"00",  X"C8",  X"FF",
  X"03",  X"01",  X"C8",  X"12",  X"4E",  X"2D",  X"18",  X"01",
  X"4E",  X"48",  X"C4",  X"0C",  X"C4",  X"30",  X"01",  X"01",
  X"02",  X"F7",  X"CC",  X"FF",  X"01",  X"2D",  X"30",  X"4C",
  X"CE",  X"00",  X"7E",  X"EC",  X"D0",  X"CC",  X"00",  X"87",
  X"00",  X"04",  X"FF",  X"01",  X"FF",  X"30",  X"FD",  X"FF",
  X"4C",  X"18",  X"2D",  X"E8",  X"97",  X"4E",  X"01",  X"00",
  X"37",  X"1C",  X"E0",  X"EA",  X"1C",  X"FA",  X"00",  X"61",
  X"EC",  X"10",  X"03",  X"02",  X"01",  X"04",  X"D4",  X"DA",
  X"D0",  X"20",  X"D0",  X"08",  X"0E",  X"D4",  X"D0",  X"14",
  X"2B",  X"11",  X"D4",  X"00",  X"29",  X"D0",  X"14",  X"18",
  X"0A",  X"A6",  X"00",  X"FF",  X"08",  X"00",  X"E0",  X"D4",
  X"1D",  X"D0",  X"EC",  X"18",  X"0A",  X"9A",  X"00",  X"D0",
  X"EC",  X"14",  X"D4",  X"0F",  X"00",  X"33",  X"01",  X"01",
  X"01",  X"E0",  X"2E",  X"01",  X"F0",  X"14",  X"D4",  X"D0",
  X"C1",  X"18",  X"D0",  X"08",  X"C4",  X"D4",  X"03",  X"00",
  X"00",  X"89",  X"11",  X"05",  X"00",  X"7A",  X"18",  X"08",
  X"14",  X"F2",  X"11",  X"00",  X"3A",  X"EC",  X"7D",  X"1C",
  X"D4",  X"D0",  X"A7",  X"18",  X"D4",  X"08",  X"AA",  X"D0",
  X"E8",  X"00",  X"40",  X"FC",  X"33",  X"F0",  X"A3",  X"E8",
  X"00",  X"0F",  X"14",  X"01",  X"7D",  X"18",  X"11",  X"D4",
  X"08",  X"00",  X"4B",  X"F4",  X"39",  X"3A",  X"01",  X"F4",
  X"F4",  X"00",  X"69",  X"01",  X"0A",  X"FF",  X"F4",  X"01",
  X"59",  X"FF",  X"05",  X"30",  X"01",  X"FF",  X"30",  X"FD",
  X"FF",  X"5B",  X"11",  X"01",  X"57",  X"00",  X"04",  X"D0",
  X"D4",  X"75",  X"18",  X"EC",  X"10",  X"0C",  X"08",  X"02",
  X"0C",  X"7B",  X"02",  X"18",  X"12",  X"4C",  X"01",  X"D0",
  X"BC",  X"08",  X"36",  X"F0",  X"01",  X"64",  X"E8",  X"F4",
  X"39",  X"06",  X"F4",  X"01",  X"00",  X"36",  X"01",  X"39",
  X"00",  X"27",  X"01",  X"39",  X"FB",  X"F0",  X"1F",  X"0C",
  X"1F",  X"01",  X"00",  X"28",  X"01",  X"BC",  X"F4",  X"F4",
  X"01",  X"B9",  X"00",  X"B1",  X"F4",  X"0F",  X"00",  X"00",
  X"A2",  X"12",  X"62",  X"00",  X"5A",  X"1C",  X"A0",  X"00",
  X"50",  X"2D",  X"0C",  X"00",  X"44",  X"00",  X"2D",  X"F0",
  X"00",  X"07",  X"0C",  X"38",  X"00",  X"3F",  X"00",  X"0C",
  X"10",  X"10",  X"08",  X"28",  X"10",  X"10",  X"00",  X"23",
  X"03",  X"00",  X"00",  X"11",  X"03",  X"00",  X"14",  X"00",
  X"08",  X"08",  X"1F",  X"00",  X"08",  X"00",  X"1A",  X"0C",
  X"24",  X"1C",  X"11",  X"00",  X"10",  X"00",  X"F6",  X"08",
  X"0C",  X"40",  X"FF",  X"00",  X"0A",  X"0C",  X"EB",  X"58",
  X"06",  X"FF",  X"10",  X"00",  X"07",  X"00",  X"08",  X"01",
  X"00",  X"FD",  X"00",  X"DE",  X"58",  X"00",  X"08",  X"01",
  X"C3",  X"58",  X"BD",  X"2D",  X"67",  X"00",  X"C2",  X"0C",
  X"28",  X"17",  X"FA",  X"58",  X"00",  X"22",  X"44",  X"00",
  X"F4",  X"00",  X"00",  X"2D",  X"28",  X"00",  X"F7",  X"00",
  X"00",  X"A0",  X"0C",  X"00",  X"04",  X"00",  X"BB",  X"58",
  X"08",  X"00",  X"30",  X"CC",  X"00",  X"B4",  X"00",  X"00",
  X"A0",  X"2D",  X"F0",  X"17",  X"D8",  X"E4",  X"F4",  X"00",
  X"00",  X"A0",  X"0C",  X"00",  X"04",  X"00",  X"8D",  X"58",
  X"08",  X"00",  X"30",  X"CC",  X"00",  X"86",  X"00",  X"00",
  X"A0",  X"F9",  X"17",  X"2D",  X"F0",  X"BF",  X"44",  X"00",
  X"90",  X"21",  X"E0",  X"20",  X"21",  X"88",  X"24",  X"21",
  X"30",  X"1C",  X"28",  X"0C",  X"0E",  X"00",  X"04",  X"08",
  X"10",  X"14",  X"18",  X"21",  X"14",  X"2C",  X"F4",  X"85",
  X"10",  X"10",  X"98",  X"01",  X"10",  X"46",  X"58",  X"88",
  X"10",  X"08",  X"00",  X"A0",  X"17",  X"B4",  X"3C",  X"01",
  X"38",  X"03",  X"04",  X"E4",  X"E0",  X"EC",  X"E8",  X"18",
  X"06",  X"CF",  X"00",  X"08",  X"18",  X"18",  X"0A",  X"C9",
  X"01",  X"0C",  X"0A",  X"C5",  X"02",  X"00",  X"A0",  X"02",
  X"04",  X"01",  X"04",  X"18",  X"01",  X"81",  X"0C",  X"00",
  X"08",  X"0C",  X"04",  X"00",  X"08",  X"10",  X"F9",  X"00",
  X"08",  X"00",  X"90",  X"9F",  X"00",  X"2D",  X"28",  X"38",
  X"00",  X"32",  X"00",  X"E0",  X"04",  X"FF",  X"06",  X"08",
  X"26",  X"00",  X"23",  X"CC",  X"0C",  X"00",  X"FC",  X"FF",
  X"FF",  X"0E",  X"01",  X"0C",  X"F4",  X"2F",  X"11",  X"01",
  X"42",  X"11",  X"11",  X"F0",  X"58",  X"32",  X"11",  X"63",
  X"00",  X"00",  X"08",  X"04",  X"10",  X"14",  X"18",  X"30",
  X"34",  X"44",  X"48",  X"08",  X"10",  X"00",  X"00",  X"08",
  X"18",  X"D3",  X"08",  X"98",  X"11",  X"CF",  X"E0",  X"AF",
  X"04",  X"00",  X"F7",  X"00",  X"46",  X"00",  X"0C",  X"EC",
  X"00",  X"A0",  X"E8",  X"18",  X"2F",  X"48",  X"08",  X"04",
  X"FC",  X"EF",  X"19",  X"00",  X"00",  X"FF",  X"09",  X"18",
  X"E0",  X"00",  X"08",  X"11",  X"01",  X"07",  X"18",  X"18",
  X"CC",  X"00",  X"08",  X"00",  X"D4",  X"19",  X"FF",  X"0E",
  X"19",  X"08",  X"01",  X"31",  X"04",  X"18",  X"01",  X"1C",
  X"19",  X"BB",  X"1C",  X"08",  X"00",  X"18",  X"C2",  X"00",
  X"08",  X"01",  X"0F",  X"E4",  X"30",  X"54",  X"03",  X"31",
  X"01",  X"1C",  X"DD",  X"04",  X"A0",  X"00",  X"50",  X"00",
  X"AA",  X"18",  X"F8",  X"04",  X"FE",  X"2F",  X"01",  X"48",
  X"04",  X"08",  X"03",  X"63",  X"FC",  X"04",  X"01",  X"0E",
  X"00",  X"F8",  X"0C",  X"0C",  X"08",  X"08",  X"0C",  X"06",
  X"01",  X"0C",  X"0C",  X"00",  X"08",  X"0D",  X"04",  X"01",
  X"0A",  X"01",  X"00",  X"2D",  X"0D",  X"08",  X"0C",  X"0C",
  X"08",  X"01",  X"01",  X"00",  X"20",  X"04",  X"FF",  X"30",
  X"03",  X"09",  X"04",  X"52",  X"5B",  X"06",  X"38",  X"03",
  X"0D",  X"08",  X"0D",  X"08",  X"04",  X"52",  X"04",  X"03",
  X"08",  X"0C",  X"04",  X"FC",  X"04",  X"FA",  X"08",  X"0C",
  X"0C",  X"08",  X"0C",  X"08",  X"58",  X"00",  X"08",  X"00",
  X"08",  X"2F",  X"50",  X"0B",  X"D3",  X"0C",  X"0C",  X"08",
  X"01",  X"08",  X"01",  X"0C",  X"04",  X"47",  X"00",  X"03",
  X"03",  X"08",  X"0C",  X"08",  X"04",  X"0C",  X"08",  X"02",
  X"01",  X"01",  X"01",  X"04",  X"38",  X"00",  X"01",  X"09",
  X"01",  X"F8",  X"0C",  X"0C",  X"08",  X"0C",  X"08",  X"0C",
  X"08",  X"01",  X"04",  X"30",  X"50",  X"02",  X"CE",  X"31",
  X"10",  X"40",  X"18",  X"21",  X"00",  X"14",  X"B2",  X"03",
  X"54",  X"0D",  X"54",  X"0C",  X"6E",  X"AB",  X"03",  X"02",
  X"01",  X"0C",  X"01",  X"04",  X"B4",  X"03",  X"06",  X"54",
  X"0F",  X"77",  X"9E",  X"03",  X"F0",  X"9B",  X"7E",  X"12",
  X"7C",  X"97",  X"03",  X"A0",  X"08",  X"00",  X"29",  X"18",
  X"0C",  X"08",  X"F3",  X"02",  X"10",  X"00",  X"F0",  X"10",
  X"02",  X"00",  X"00",  X"1F",  X"00",  X"00",  X"15",  X"13",
  X"00",  X"03",  X"12",  X"00",  X"24",  X"00",  X"1C",  X"00",
  X"98",  X"08",  X"08",  X"08",  X"00",  X"0A",  X"08",  X"08",
  X"00",  X"EF",  X"13",  X"00",  X"04",  X"E8",  X"08",  X"00",
  X"08",  X"00",  X"2D",  X"01",  X"F0",  X"4E",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"2B",  X"00",  X"00",  X"B5",  X"16",
  X"13",  X"03",  X"14",  X"13",  X"14",  X"08",  X"12",  X"12",
  X"8D",  X"00",  X"10",  X"01",  X"8A",  X"0A",  X"16",  X"2C",
  X"12",  X"00",  X"12",  X"00",  X"A2",  X"10",  X"00",  X"62",
  X"0C",  X"12",  X"88",  X"00",  X"08",  X"12",  X"00",  X"D0",
  X"08",  X"12",  X"00",  X"DA",  X"12",  X"00",  X"04",  X"00",
  X"D2",  X"08",  X"00",  X"15",  X"05",  X"15",  X"12",  X"12",
  X"15",  X"0A",  X"14",  X"08",  X"00",  X"13",  X"15",  X"08",
  X"00",  X"12",  X"12",  X"08",  X"13",  X"00",  X"B1",  X"08",
  X"0C",  X"15",  X"15",  X"00",  X"1E",  X"00",  X"10",  X"10",
  X"00",  X"1C",  X"08",  X"13",  X"DE",  X"13",  X"80",  X"DC",
  X"00",  X"10",  X"00",  X"00",  X"09",  X"15",  X"0C",  X"13",
  X"00",  X"6D",  X"15",  X"14",  X"10",  X"00",  X"08",  X"12",
  X"CB",  X"12",  X"04",  X"E0",  X"08",  X"12",  X"00",  X"16",
  X"13",  X"10",  X"01",  X"13",  X"14",  X"14",  X"CD",  X"13",
  X"00",  X"13",  X"00",  X"43",  X"10",  X"00",  X"C6",  X"08",
  X"0C",  X"40",  X"0C",  X"08",  X"FF",  X"14",  X"0A",  X"0B",
  X"14",  X"24",  X"1C",  X"00",  X"14",  X"00",  X"F3",  X"0C",
  X"B3",  X"13",  X"B1",  X"12",  X"08",  X"00",  X"12",  X"12",
  X"08",  X"00",  X"12",  X"A8",  X"12",  X"0A",  X"13",  X"16",
  X"24",  X"1C",  X"00",  X"16",  X"00",  X"DC",  X"0C",  X"12",
  X"7D",  X"08",  X"14",  X"10",  X"00",  X"D3",  X"00",  X"76",
  X"08",  X"92",  X"15",  X"08",  X"00",  X"15",  X"15",  X"08",
  X"00",  X"68",  X"15",  X"0A",  X"13",  X"0B",  X"01",  X"00",
  X"48",  X"01",  X"01",  X"45",  X"16",  X"10",  X"64",  X"FF",
  X"00",  X"2F",  X"00",  X"0C",  X"0C",  X"01",  X"00",  X"55",
  X"10",  X"B0",  X"0C",  X"A0",  X"6E",  X"18",  X"E0",  X"31",
  X"00",  X"04",  X"FF",  X"14",  X"08",  X"28",  X"00",  X"0E",
  X"11",  X"FF",  X"06",  X"10",  X"00",  X"00",  X"0C",  X"08",
  X"00",  X"16",  X"58",  X"FF",  X"19",  X"00",  X"CC",  X"0C",
  X"10",  X"00",  X"FA",  X"FF",  X"10",  X"00",  X"EA",  X"0E",
  X"58",  X"D2",  X"14",  X"0C",  X"00",  X"E2",  X"0C",  X"E2",
  X"14",  X"FF",  X"ED",  X"CC",  X"00",  X"00",  X"D4",  X"04",
  X"22",  X"00",  X"08",  X"00",  X"A0",  X"35",  X"00",  X"E0",
  X"30",  X"00",  X"04",  X"FF",  X"13",  X"08",  X"27",  X"00",
  X"0E",  X"FF",  X"06",  X"10",  X"00",  X"00",  X"0C",  X"08",
  X"00",  X"16",  X"58",  X"FF",  X"19",  X"00",  X"CC",  X"0C",
  X"10",  X"00",  X"FA",  X"FF",  X"10",  X"00",  X"EB",  X"0E",
  X"58",  X"9A",  X"13",  X"0C",  X"00",  X"E3",  X"0C",  X"AA",
  X"13",  X"FF",  X"ED",  X"CC",  X"00",  X"00",  X"D5",  X"04",
  X"EA",  X"00",  X"08",  X"00",  X"2D",  X"08",  X"78",  X"2D",
  X"08",  X"48",  X"2D",  X"08",  X"48",  X"A0",  X"18",  X"00",
  X"2D",  X"14",  X"30",  X"1A",  X"18",  X"1F",  X"2D",  X"00",
  X"06",  X"1A",  X"34",  X"30",  X"08",  X"30",  X"2D",  X"00",
  X"14",  X"48",  X"00",  X"F8",  X"34",  X"08",  X"00",  X"08",
  X"2D",  X"F0",  X"09",  X"01",  X"00",  X"E0",  X"00",  X"00",
  X"60",  X"0C",  X"02",  X"3B",  X"43",  X"0E",  X"00",  X"17",
  X"2D",  X"F0",  X"06",  X"C0",  X"00",  X"10",  X"C8",  X"3C",
  X"01",  X"08",  X"02",  X"02",  X"20",  X"FF",  X"02",  X"2D",
  X"28",  X"0C",  X"00",  X"06",  X"0C",  X"0C",  X"00",  X"00",
  X"0C",  X"F0",  X"84",  X"00",  X"00",  X"29",  X"2D",  X"0C",
  X"F0",  X"80",  X"10",  X"00",  X"0C",  X"17",  X"B4",  X"3C",
  X"00",  X"00",  X"0A",  X"14",  X"AA",  X"0E",  X"00",  X"1F",
  X"00",  X"0C",  X"01",  X"0C",  X"08",  X"00",  X"10",  X"00",
  X"01",  X"14",  X"08",  X"00",  X"21",  X"30",  X"01",  X"D3",
  X"0C",  X"00",  X"00",  X"4C",  X"D5",  X"0C",  X"0C",  X"02",
  X"43",  X"10",  X"00",  X"0C",  X"01",  X"14",  X"08",  X"00",
  X"A0",  X"FF",  X"03",  X"29",  X"18",  X"03",  X"2E",  X"08",
  X"BF",  X"19",  X"20",  X"08",  X"FF",  X"19",  X"80",  X"08",
  X"19",  X"00",  X"01",  X"04",  X"01",  X"03",  X"12",  X"FC",
  X"00",  X"19",  X"20",  X"00",  X"01",  X"19",  X"1A",  X"01",
  X"02",  X"19",  X"16",  X"02",  X"03",  X"19",  X"12",  X"03",
  X"03",  X"E8",  X"04",  X"18",  X"00",  X"08",  X"00",  X"08",
  X"00",  X"00",  X"FD",  X"01",  X"00",  X"19",  X"FB",  X"FF",
  X"08",  X"01",  X"08",  X"00",  X"A0",  X"0F",  X"18",  X"19",
  X"06",  X"1A",  X"18",  X"03",  X"0D",  X"19",  X"00",  X"08",
  X"00",  X"01",  X"01",  X"01",  X"03",  X"FD",  X"01",  X"08",
  X"00",  X"18",  X"00",  X"00",  X"F0",  X"0F",  X"04",  X"04",
  X"08",  X"08",  X"0C",  X"0C",  X"10",  X"F5",  X"10",  X"F0",
  X"04",  X"04",  X"01",  X"01",  X"04",  X"03",  X"0D",  X"1A",
  X"DE",  X"0D",  X"00",  X"01",  X"01",  X"04",  X"01",  X"03",
  X"FC",  X"01",  X"FC",  X"02",  X"02",  X"01",  X"03",  X"02",
  X"01",  X"CD",  X"01",  X"A0",  X"19",  X"18",  X"19",  X"13",
  X"1A",  X"1A",  X"01",  X"10",  X"0F",  X"00",  X"0A",  X"FF",
  X"1A",  X"FF",  X"00",  X"FF",  X"FF",  X"FF",  X"FB",  X"00",
  X"08",  X"00",  X"0F",  X"0D",  X"18",  X"00",  X"FA",  X"00",
  X"01",  X"01",  X"01",  X"03",  X"FD",  X"01",  X"08",  X"00",
  X"03",  X"F5",  X"00",  X"1A",  X"19",  X"18",  X"00",  X"00",
  X"F0",  X"0F",  X"04",  X"04",  X"08",  X"08",  X"0C",  X"0C",
  X"10",  X"F5",  X"10",  X"F0",  X"04",  X"04",  X"01",  X"01",
  X"04",  X"03",  X"0D",  X"1A",  X"D9",  X"0D",  X"00",  X"01",
  X"01",  X"04",  X"01",  X"03",  X"FC",  X"01",  X"FC",  X"02",
  X"02",  X"01",  X"03",  X"02",  X"01",  X"C8",  X"01",  X"A0",
  X"FF",  X"03",  X"2A",  X"18",  X"03",  X"2A",  X"00",  X"08",
  X"03",  X"0F",  X"10",  X"18",  X"01",  X"1A",  X"11",  X"18",
  X"00",  X"04",  X"08",  X"0C",  X"F0",  X"0F",  X"FA",  X"10",
  X"F0",  X"0F",  X"F0",  X"03",  X"10",  X"0E",  X"0D",  X"00",
  X"01",  X"04",  X"01",  X"03",  X"FD",  X"01",  X"FC",  X"03",
  X"FC",  X"04",  X"01",  X"0D",  X"00",  X"07",  X"00",  X"01",
  X"01",  X"1A",  X"FE",  X"01",  X"08",  X"00",  X"00",  X"08",
  X"00",  X"4C",  X"04",  X"02",  X"01",  X"00",  X"01",  X"08",
  X"00",  X"08",  X"C0",  X"02",  X"04",  X"00",  X"10",  X"10",
  X"00",  X"02",  X"04",  X"00",  X"08",  X"08",  X"02",  X"04",
  X"00",  X"04",  X"04",  X"02",  X"05",  X"00",  X"02",  X"02",
  X"00",  X"05",  X"00",  X"02",  X"04",  X"01",  X"08",  X"00",
  X"08",  X"20",  X"00",  X"07",  X"0C",  X"3F",  X"01",  X"07",
  X"00",  X"02",  X"2C",  X"02",  X"02",  X"00",  X"08",  X"02",
  X"FF",  X"02",  X"1B",  X"00",  X"FF",  X"05",  X"0F",  X"08",
  X"08",  X"0F",  X"05",  X"03",  X"04",  X"04",  X"03",  X"05",
  X"01",  X"02",  X"02",  X"01",  X"07",  X"00",  X"01",  X"00",
  X"0B",  X"01",  X"00",  X"08",  X"02",  X"10",  X"FF",  X"EA",
  X"10",  X"E7",  X"08",  X"20",  X"08",  X"02",  X"01",  X"01",
  X"00",  X"08",  X"02",  X"A0",  X"18",  X"10",  X"10",  X"02",
  X"11",  X"04",  X"02",  X"02",  X"02",  X"04",  X"04",  X"14",
  X"FC",  X"FC",  X"00",  X"00",  X"04",  X"06",  X"02",  X"FA",
  X"FC",  X"08",  X"00",  X"04",  X"00",  X"01",  X"08",  X"00",
  X"00",  X"00",  X"01",  X"02",  X"00",  X"08",  X"98",  X"01",
  X"00",  X"60",  X"60",  X"08",  X"98",  X"01",  X"14",  X"13",
  X"11",  X"00",  X"EC",  X"1E",  X"08",  X"01",  X"00",  X"04",
  X"60",  X"60",  X"08",  X"98",  X"01",  X"00",  X"01",  X"F9",
  X"04",  X"00",  X"01",  X"60",  X"60",  X"08",  X"98",  X"98",
  X"10",  X"04",  X"02",  X"10",  X"5D",  X"11",  X"20",  X"08",
  X"00",  X"10",  X"0A",  X"13",  X"14",  X"0B",  X"10",  X"08",
  X"04",  X"00",  X"FC",  X"02",  X"02",  X"15",  X"00",  X"08",
  X"04",  X"11",  X"F8",  X"F8",  X"08",  X"00",  X"10",  X"1E",
  X"00",  X"F5",  X"15",  X"00",  X"20",  X"18",  X"08",  X"04",
  X"00",  X"FC",  X"02",  X"08",  X"02",  X"00",  X"08",  X"0D",
  X"02",  X"01",  X"F8",  X"F8",  X"08",  X"00",  X"00",  X"01",
  X"04",  X"F8",  X"F8",  X"08",  X"00",  X"FC",  X"F5",  X"F7",
  X"FC",  X"E4",  X"20",  X"88",  X"FC",  X"BA",  X"18",  X"20",
  X"F8",  X"19",  X"F0",  X"B4",  X"F4",  X"10",  X"10",  X"F8",
  X"FC",  X"01",  X"02",  X"F4",  X"05",  X"F0",  X"02",  X"00",
  X"0C",  X"20",  X"EC",  X"14",  X"EC",  X"02",  X"EC",  X"EC",
  X"2A",  X"C0",  X"08",  X"00",  X"EC",  X"14",  X"EC",  X"01",
  X"EC",  X"EC",  X"2C",  X"C0",  X"08",  X"00",  X"17",  X"0A",
  X"2D",  X"10",  X"2D",  X"18",  X"FF",  X"FF",  X"48",  X"08",
  X"00",  X"03",  X"2D",  X"80",  X"08",  X"08",  X"A0",  X"4C",
  X"00",  X"0D",  X"18",  X"02",  X"02",  X"00",  X"13",  X"10",
  X"00",  X"02",  X"10",  X"0C",  X"08",  X"00",  X"18",  X"04",
  X"DD",  X"10",  X"4C",  X"08",  X"00",  X"EE",  X"00",  X"08",
  X"00",  X"01",  X"01",  X"19",  X"05",  X"D0",  X"02",  X"00",
  X"F7",  X"00",  X"04",  X"08",  X"10",  X"0C",  X"08",  X"00",
  X"90",  X"01",  X"18",  X"F0",  X"D2",  X"F4",  X"00",  X"02",
  X"F8",  X"00",  X"1A",  X"03",  X"14",  X"00",  X"05",  X"08",
  X"00",  X"03",  X"F8",  X"00",  X"1E",  X"00",  X"FC",  X"C3",
  X"FC",  X"00",  X"2A",  X"F8",  X"FC",  X"14",  X"F8",  X"01",
  X"18",  X"00",  X"01",  X"00",  X"18",  X"10",  X"CE",  X"03",
  X"00",  X"02",  X"01",  X"8E",  X"04",  X"05",  X"08",  X"00",
  X"08",  X"00",  X"A8",  X"F8",  X"F8",  X"14",  X"01",  X"10",
  X"20",  X"00",  X"EC",  X"01",  X"CD",  X"08",  X"00",  X"35",
  X"08",  X"00",  X"08",  X"00",  X"FC",  X"08",  X"02",  X"03",
  X"14",  X"08",  X"D5",  X"F8",  X"A0",  X"10",  X"10",  X"01",
  X"4A",  X"18",  X"00",  X"61",  X"19",  X"00",  X"14",  X"7F",
  X"04",  X"10",  X"10",  X"04",  X"0C",  X"02",  X"04",  X"01",
  X"02",  X"3F",  X"09",  X"04",  X"04",  X"FF",  X"14",  X"14",
  X"00",  X"00",  X"00",  X"10",  X"0C",  X"10",  X"0C",  X"0B",
  X"0D",  X"02",  X"10",  X"0D",  X"02",  X"04",  X"00",  X"04",
  X"04",  X"1A",  X"EF",  X"10",  X"19",  X"12",  X"FC",  X"3F",
  X"FF",  X"00",  X"10",  X"0C",  X"03",  X"10",  X"0D",  X"02",
  X"04",  X"00",  X"10",  X"04",  X"F5",  X"10",  X"FC",  X"00",
  X"07",  X"FC",  X"FC",  X"00",  X"00",  X"FD",  X"FF",  X"10",
  X"08",  X"08",  X"04",  X"14",  X"02",  X"01",  X"01",  X"04",
  X"04",  X"FC",  X"FC",  X"00",  X"00",  X"03",  X"0B",  X"01",
  X"FA",  X"FC",  X"2C",  X"00",  X"01",  X"14",  X"10",  X"08",
  X"08",  X"03",  X"A5",  X"19",  X"01",  X"1A",  X"01",  X"A0",
  X"14",  X"A0",  X"10",  X"08",  X"01",  X"05",  X"18",  X"11",
  X"01",  X"06",  X"04",  X"01",  X"01",  X"FE",  X"01",  X"0F",
  X"12",  X"00",  X"0C",  X"14",  X"00",  X"00",  X"01",  X"11",
  X"FD",  X"04",  X"04",  X"02",  X"01",  X"04",  X"10",  X"04",
  X"1F",  X"02",  X"14",  X"04",  X"1C",  X"04",  X"20",  X"00",
  X"1A",  X"00",  X"1A",  X"0D",  X"00",  X"04",  X"00",  X"04",
  X"02",  X"F8",  X"0C",  X"00",  X"03",  X"10",  X"4C",  X"04",
  X"02",  X"01",  X"00",  X"FF",  X"01",  X"10",  X"08",  X"08",
  X"00",  X"00",  X"04",  X"02",  X"F2",  X"04",  X"00",  X"00",
  X"04",  X"02",  X"F6",  X"04",  X"EB",  X"4C",  X"98",  X"10",
  X"10",  X"11",  X"80",  X"18",  X"11",  X"10",  X"01",  X"08",
  X"11",  X"01",  X"03",  X"04",  X"01",  X"C1",  X"04",  X"14",
  X"02",  X"17",  X"04",  X"17",  X"08",  X"08",  X"1B",  X"00",
  X"04",  X"01",  X"FE",  X"00",  X"04",  X"02",  X"15",  X"14",
  X"F8",  X"04",  X"14",  X"02",  X"1C",  X"04",  X"1C",  X"47",
  X"04",  X"3F",  X"FF",  X"00",  X"11",  X"1D",  X"FC",  X"F8",
  X"1B",  X"00",  X"00",  X"FC",  X"59",  X"11",  X"00",  X"FC",
  X"11",  X"12",  X"53",  X"10",  X"19",  X"10",  X"10",  X"13",
  X"01",  X"02",  X"04",  X"00",  X"1A",  X"04",  X"EC",  X"10",
  X"00",  X"00",  X"10",  X"00",  X"1E",  X"FC",  X"00",  X"F8",
  X"19",  X"1B",  X"00",  X"00",  X"FC",  X"11",  X"37",  X"10",
  X"08",  X"12",  X"02",  X"FC",  X"00",  X"10",  X"2F",  X"10",
  X"04",  X"00",  X"04",  X"11",  X"1A",  X"19",  X"13",  X"EC",
  X"10",  X"00",  X"04",  X"1D",  X"BF",  X"04",  X"00",  X"11",
  X"10",  X"FC",  X"00",  X"09",  X"FC",  X"10",  X"08",  X"00",
  X"00",  X"00",  X"06",  X"10",  X"FF",  X"FB",  X"FC",  X"10",
  X"08",  X"00",  X"19",  X"1A",  X"83",  X"01",  X"A0",  X"01",
  X"46",  X"18",  X"01",  X"14",  X"10",  X"08",  X"08",  X"A0",
  X"10",  X"3F",  X"14",  X"FF",  X"00",  X"00",  X"15",  X"F6",
  X"1A",  X"10",  X"08",  X"F2",  X"1A",  X"10",  X"15",  X"08",
  X"10",  X"13",  X"00",  X"01",  X"04",  X"12",  X"EF",  X"10",
  X"00",  X"0C",  X"00",  X"08",  X"01",  X"0A",  X"04",  X"04",
  X"02",  X"01",  X"01",  X"10",  X"04",  X"08",  X"19",  X"01",
  X"16",  X"18",  X"10",  X"08",  X"0C",  X"02",  X"0C",  X"1D",
  X"02",  X"4C",  X"04",  X"02",  X"01",  X"00",  X"01",  X"E8",
  X"1A",  X"A0",  X"03",  X"32",  X"18",  X"02",  X"00",  X"25",
  X"00",  X"48",  X"00",  X"35",  X"10",  X"01",  X"0F",  X"19",
  X"01",  X"00",  X"1A",  X"00",  X"00",  X"00",  X"18",  X"11",
  X"08",  X"01",  X"F7",  X"01",  X"19",  X"11",  X"18",  X"10",
  X"00",  X"08",  X"01",  X"4C",  X"04",  X"02",  X"01",  X"00",
  X"01",  X"00",  X"EA",  X"08",  X"08",  X"19",  X"11",  X"07",
  X"10",  X"00",  X"00",  X"E6",  X"08",  X"FF",  X"2D",  X"02",
  X"98",  X"01",  X"19",  X"18",  X"8B",  X"00",  X"C7",  X"08",
  X"7E",  X"71",  X"48",  X"08",  X"C9",  X"00",  X"A0",  X"09",
  X"B9",  X"08",  X"18",  X"01",  X"01",  X"06",  X"00",  X"01",
  X"01",  X"FE",  X"01",  X"B3",  X"10",  X"01",  X"14",  X"10",
  X"09",  X"0A",  X"10",  X"09",  X"09",  X"11",  X"08",  X"D0",
  X"10",  X"66",  X"0A",  X"01",  X"11",  X"F9",  X"11",  X"1A",
  X"1A",  X"F8",  X"11",  X"0D",  X"00",  X"1A",  X"08",  X"D0",
  X"10",  X"56",  X"0A",  X"01",  X"11",  X"01",  X"F8",  X"1A",
  X"08",  X"08",  X"A0",  X"00",  X"04",  X"18",  X"A8",  X"1A",
  X"62",  X"18",  X"F8",  X"04",  X"0B",  X"16",  X"09",  X"02",
  X"10",  X"00",  X"1A",  X"09",  X"10",  X"08",  X"00",  X"F8",
  X"11",  X"1A",  X"FB",  X"1F",  X"FF",  X"F8",  X"FC",  X"03",
  X"54",  X"17",  X"2F",  X"48",  X"08",  X"17",  X"01",  X"F5",
  X"10",  X"04",  X"FE",  X"0D",  X"04",  X"01",  X"64",  X"00",
  X"FC",  X"17",  X"03",  X"61",  X"08",  X"01",  X"A0",  X"00",
  X"F8",  X"13",  X"04",  X"F8",  X"FC",  X"04",  X"5D",  X"17",
  X"02",  X"03",  X"C9",  X"08",  X"02",  X"03",  X"91",  X"1A",
  X"0C",  X"08",  X"FC",  X"08",  X"08",  X"24",  X"C8",  X"0C",
  X"13",  X"19",  X"18",  X"08",  X"00",  X"08",  X"1B",  X"10",
  X"04",  X"0C",  X"10",  X"08",  X"08",  X"10",  X"24",  X"18",
  X"04",  X"14",  X"08",  X"08",  X"00",  X"18",  X"20",  X"04",
  X"1C",  X"08",  X"00",  X"00",  X"08",  X"13",  X"04",  X"04",
  X"08",  X"08",  X"04",  X"04",  X"16",  X"08",  X"11",  X"0F",
  X"0D",  X"11",  X"01",  X"12",  X"04",  X"12",  X"04",  X"01",
  X"04",  X"E3",  X"10",  X"08",  X"00",  X"01",  X"11",  X"04",
  X"01",  X"04",  X"03",  X"10",  X"04",  X"01",  X"04",  X"2D",
  X"08",  X"F0",  X"A3",  X"00",  X"0C",  X"08",  X"02",  X"0C",
  X"16",  X"DD",  X"08",  X"17",  X"10",  X"12",  X"01",  X"A7",
  X"03",  X"0C",  X"08",  X"FC",  X"08",  X"08",  X"24",  X"94",
  X"0C",  X"13",  X"19",  X"18",  X"18",  X"00",  X"08",  X"1B",
  X"10",  X"04",  X"0C",  X"10",  X"08",  X"08",  X"10",  X"24",
  X"18",  X"04",  X"14",  X"08",  X"08",  X"00",  X"18",  X"20",
  X"04",  X"1C",  X"08",  X"00",  X"00",  X"04",  X"04",  X"08",
  X"08",  X"11",  X"11",  X"01",  X"04",  X"08",  X"10",  X"04",
  X"01",  X"01",  X"92",  X"04",  X"08",  X"00",  X"1A",  X"D7",
  X"10",  X"00",  X"2D",  X"F8",  X"04",  X"FE",  X"03",  X"03",
  X"55",  X"FC",  X"24",  X"4C",  X"13",  X"19",  X"18",  X"18",
  X"00",  X"00",  X"1B",  X"08",  X"04",  X"04",  X"10",  X"08",
  X"08",  X"08",  X"24",  X"10",  X"0C",  X"0C",  X"08",  X"10",
  X"10",  X"10",  X"18",  X"18",  X"14",  X"14",  X"00",  X"00",
  X"04",  X"04",  X"08",  X"08",  X"19",  X"B7",  X"10",  X"5D",
  X"10",  X"08",  X"00",  X"0C",  X"FC",  X"08",  X"0C",  X"08",
  X"24",  X"0C",  X"08",  X"08",  X"3C",  X"0C",  X"19",  X"85",
  X"08",  X"13",  X"5C",  X"04",  X"04",  X"FC",  X"17",  X"01",
  X"15",  X"04",  X"11",  X"11",  X"01",  X"04",  X"08",  X"10",
  X"04",  X"01",  X"01",  X"39",  X"04",  X"08",  X"19",  X"6D",
  X"19",  X"D4",  X"19",  X"12",  X"17",  X"04",  X"FC",  X"16",
  X"17",  X"3D",  X"08",  X"19",  X"60",  X"18",  X"8C",  X"11",
  X"A0",  X"00",  X"1F",  X"2D",  X"48",  X"00",  X"14",  X"3C",
  X"04",  X"FF",  X"0C",  X"00",  X"01",  X"02",  X"11",  X"00",
  X"00",  X"FC",  X"FF",  X"FD",  X"00",  X"00",  X"00",  X"F2",
  X"04",  X"3C",  X"00",  X"04",  X"00",  X"00",  X"18",  X"08",
  X"00",  X"E3",  X"F0",  X"A0",  X"00",  X"00",  X"04",  X"00",
  X"FB",  X"18",  X"52",  X"00",  X"00",  X"A0",  X"2D",  X"F0",
  X"01",  X"32",  X"00",  X"4C",  X"00",  X"16",  X"48",  X"00",
  X"11",  X"00",  X"0B",  X"04",  X"10",  X"18",  X"3E",  X"00",
  X"00",  X"FC",  X"10",  X"4C",  X"04",  X"3C",  X"F3",  X"11",
  X"34",  X"18",  X"48",  X"00",  X"0E",  X"54",  X"4C",  X"11",
  X"0A",  X"54",  X"10",  X"18",  X"28",  X"00",  X"10",  X"FC",
  X"10",  X"54",  X"00",  X"05",  X"38",  X"1F",  X"18",  X"38",
  X"00",  X"04",  X"3C",  X"08",  X"00",  X"00",  X"18",  X"E0",
  X"00",  X"FA",  X"00",  X"B8",  X"00",  X"00",  X"09",  X"00",
  X"09",  X"00",  X"1F",  X"04",  X"04",  X"01",  X"01",  X"01",
  X"1F",  X"08",  X"01",  X"00",  X"01",  X"09",  X"09",  X"1F",
  X"01",  X"00",  X"08",  X"08",  X"1F",  X"0E",  X"2D",  X"F0",
  X"00",  X"DC",  X"00",  X"00",  X"A0",  X"2D",  X"0E",  X"F0",
  X"19",  X"58",  X"1A",  X"FF",  X"08",  X"04",  X"0C",  X"01",
  X"50",  X"0C",  X"08",  X"08",  X"0C",  X"04",  X"02",  X"0C",
  X"08",  X"08",  X"A0",  X"0C",  X"18",  X"00",  X"19",  X"1A",
  X"08",  X"2D",  X"F0",  X"0E",  X"00",  X"3C",  X"02",  X"0C",
  X"04",  X"02",  X"F0",  X"0E",  X"0C",  X"76",  X"11",  X"00",
  X"A0",  X"2D",  X"0E",  X"F0",  X"19",  X"3E",  X"1A",  X"00",
  X"07",  X"0C",  X"50",  X"08",  X"50",  X"08",  X"08",  X"04",
  X"02",  X"0C",  X"08",  X"08",  X"08",  X"03",  X"1E",  X"00",
  X"00",  X"00",  X"02",  X"18",  X"BF",  X"20",  X"FF",  X"80",
  X"02",  X"02",  X"01",  X"03",  X"09",  X"04",  X"08",  X"00",
  X"01",  X"03",  X"22",  X"00",  X"04",  X"04",  X"00",  X"00",
  X"02",  X"F7",  X"04",  X"00",  X"00",  X"0A",  X"00",  X"11",
  X"00",  X"01",  X"00",  X"01",  X"00",  X"0A",  X"00",  X"00",
  X"02",  X"F8",  X"00",  X"FF",  X"FF",  X"08",  X"01",  X"00",
  X"FF",  X"FF",  X"08",  X"01",  X"08",  X"00",  X"A0",  X"03",
  X"1C",  X"18",  X"00",  X"BF",  X"FF",  X"0D",  X"01",  X"20",
  X"80",  X"04",  X"12",  X"18",  X"04",  X"00",  X"0D",  X"02",
  X"04",  X"0C",  X"00",  X"04",  X"00",  X"0D",  X"02",  X"04",
  X"F5",  X"04",  X"03",  X"00",  X"00",  X"00",  X"FE",  X"01",
  X"18",  X"08",  X"00",  X"A0",  X"32",  X"19",  X"1A",  X"80",
  X"A5",  X"1B",  X"FF",  X"04",  X"80",  X"08",  X"08",  X"00",
  X"FD",  X"00",  X"00",  X"08",  X"08",  X"A0",  X"19",  X"CE",
  X"1A",  X"08",  X"2C",  X"18",  X"00",  X"1E",  X"00",  X"FC",
  X"FC",  X"FC",  X"24",  X"16",  X"13",  X"0F",  X"18",  X"00",
  X"04",  X"1B",  X"0A",  X"08",  X"08",  X"0C",  X"24",  X"05",
  X"10",  X"10",  X"14",  X"18",  X"08",  X"00",  X"04",  X"08",
  X"00",  X"8E",  X"00",  X"08",  X"00",  X"A0",  X"32",  X"19",
  X"37",  X"80",  X"FF",  X"04",  X"80",  X"08",  X"08",  X"00",
  X"FD",  X"00",  X"00",  X"08",  X"08",  X"A0",  X"00",  X"3E",
  X"00",  X"21",  X"58",  X"0C",  X"00",  X"3A",  X"00",  X"2D",
  X"F0",  X"00",  X"07",  X"0C",  X"38",  X"00",  X"3B",  X"00",
  X"0C",  X"10",  X"00",  X"30",  X"10",  X"08",  X"3F",  X"00",
  X"2C",  X"00",  X"08",  X"0C",  X"00",  X"1C",  X"00",  X"02",
  X"FF",  X"0C",  X"80",  X"2E",  X"10",  X"30",  X"00",  X"08",
  X"40",  X"01",  X"05",  X"30",  X"D8",  X"F0",  X"30",  X"44",
  X"00",  X"06",  X"0C",  X"D1",  X"F0",  X"44",  X"0C",  X"8A",
  X"12",  X"67",  X"12",  X"CF",  X"00",  X"08",  X"10",  X"6C",
  X"12",  X"C7",  X"2D",  X"7E",  X"12",  X"C5",  X"00",  X"08",
  X"10",  X"0A",  X"00",  X"0C",  X"10",  X"00",  X"C7",  X"10",
  X"F3",  X"B3",  X"18",  X"D3",  X"30",  X"49",  X"19",  X"C1",
  X"08",  X"08",  X"2D",  X"F0",  X"00",  X"A0",  X"00",  X"00",
  X"A0",  X"32",  X"19",  X"1A",  X"C5",  X"80",  X"FF",  X"04",
  X"80",  X"08",  X"08",  X"00",  X"FD",  X"00",  X"00",  X"08",
  X"08",  X"A0",  X"32",  X"19",  X"1A",  X"80",  X"BA",  X"1B",
  X"FF",  X"04",  X"80",  X"08",  X"08",  X"00",  X"FD",  X"00",
  X"00",  X"08",  X"08",  X"A0",  X"32",  X"19",  X"1A",  X"80",
  X"AF",  X"1B",  X"FF",  X"04",  X"80",  X"08",  X"08",  X"00",
  X"FD",  X"00",  X"00",  X"08",  X"08",  X"09",  X"00",  X"FF",
  X"25",  X"00",  X"09",  X"09",  X"09",  X"09",  X"09",  X"09",
  X"09",  X"09",  X"09",  X"09",  X"09",  X"09",  X"09",  X"09",
  X"09",  X"09",  X"09",  X"09",  X"09",  X"09",  X"09",  X"09",
  X"09",  X"09",  X"09",  X"09",  X"09",  X"09",  X"09",  X"09",
  X"09",  X"09",  X"00",  X"08",  X"00",  X"09",  X"09",  X"09",
  X"09",  X"09",  X"09",  X"09",  X"09",  X"09",  X"09",  X"09",
  X"09",  X"00",  X"00",  X"0C",  X"14",  X"08",  X"0C",  X"0B",
  X"00",  X"08",  X"08",  X"08",  X"00",  X"04",  X"00",  X"03",
  X"09",  X"08",  X"00",  X"05",  X"08",  X"02",  X"08",  X"00",
  X"0D",  X"95",  X"00",  X"00",  X"01",  X"28",  X"00",  X"01",
  X"0D",  X"01",  X"04",  X"FC",  X"01",  X"0D",  X"07",  X"01",
  X"04",  X"01",  X"01",  X"07",  X"01",  X"0B",  X"F7",  X"00",
  X"02",  X"00",  X"01",  X"76",  X"00",  X"0D",  X"01",  X"0A",
  X"00",  X"01",  X"05",  X"01",  X"0D",  X"04",  X"01",  X"0D",
  X"01",  X"01",  X"F7",  X"00",  X"65",  X"04",  X"0B",  X"FE",
  X"01",  X"65",  X"01",  X"00",  X"04",  X"2F",  X"01",  X"0D",
  X"17",  X"01",  X"0D",  X"0B",  X"01",  X"0D",  X"05",  X"01",
  X"0D",  X"50",  X"0F",  X"0D",  X"4D",  X"0D",  X"0D",  X"05",
  X"01",  X"0D",  X"47",  X"0B",  X"0D",  X"44",  X"09",  X"0D",
  X"0B",  X"01",  X"0D",  X"05",  X"01",  X"0D",  X"3B",  X"07",
  X"0D",  X"38",  X"05",  X"0D",  X"05",  X"01",  X"0D",  X"32",
  X"03",  X"0D",  X"2F",  X"01",  X"0D",  X"17",  X"01",  X"0D",
  X"0B",  X"01",  X"0D",  X"05",  X"01",  X"0D",  X"23",  X"FF",
  X"0D",  X"20",  X"FD",  X"0D",  X"05",  X"01",  X"0D",  X"1A",
  X"FB",  X"0D",  X"17",  X"F9",  X"0D",  X"0B",  X"01",  X"0D",
  X"05",  X"01",  X"0D",  X"0E",  X"F7",  X"0D",  X"0B",  X"F5",
  X"0D",  X"05",  X"01",  X"0D",  X"05",  X"F3",  X"0D",  X"02",
  X"F1",  X"01",  X"A2",  X"00",  X"02",  X"01",  X"00",  X"02",
  X"0A",  X"08",  X"0A",  X"0B",  X"00",  X"08",  X"08",  X"08",
  X"00",  X"04",  X"00",  X"03",  X"09",  X"08",  X"00",  X"05",
  X"08",  X"02",  X"08",  X"00",  X"0D",  X"95",  X"00",  X"00",
  X"01",  X"28",  X"00",  X"01",  X"0D",  X"01",  X"04",  X"FC",
  X"01",  X"0D",  X"07",  X"01",  X"04",  X"01",  X"01",  X"07",
  X"01",  X"0B",  X"F7",  X"00",  X"02",  X"00",  X"01",  X"76",
  X"00",  X"0D",  X"01",  X"0A",  X"00",  X"01",  X"05",  X"01",
  X"0D",  X"04",  X"01",  X"0D",  X"01",  X"01",  X"F7",  X"00",
  X"65",  X"04",  X"0B",  X"FE",  X"01",  X"65",  X"01",  X"00",
  X"04",  X"2F",  X"01",  X"0D",  X"17",  X"01",  X"0D",  X"0B",
  X"01",  X"0D",  X"05",  X"01",  X"0D",  X"50",  X"0F",  X"0D",
  X"4D",  X"0D",  X"0D",  X"05",  X"01",  X"0D",  X"47",  X"0B",
  X"0D",  X"44",  X"09",  X"0D",  X"0B",  X"01",  X"0D",  X"05",
  X"01",  X"0D",  X"3B",  X"07",  X"0D",  X"38",  X"05",  X"0D",
  X"05",  X"01",  X"0D",  X"32",  X"03",  X"0D",  X"2F",  X"01",
  X"0D",  X"17",  X"01",  X"0D",  X"0B",  X"01",  X"0D",  X"05",
  X"01",  X"0D",  X"23",  X"FF",  X"0D",  X"20",  X"FD",  X"0D",
  X"05",  X"01",  X"0D",  X"1A",  X"FB",  X"0D",  X"17",  X"F9",
  X"0D",  X"0B",  X"01",  X"0D",  X"05",  X"01",  X"0D",  X"0E",
  X"F7",  X"0D",  X"0B",  X"F5",  X"0D",  X"05",  X"01",  X"0D",
  X"05",  X"F3",  X"0D",  X"02",  X"F1",  X"01",  X"A2",  X"00",
  X"02",  X"09",  X"00",  X"02",  X"0B",  X"08",  X"0B",  X"08",
  X"00",  X"08",  X"00",  X"08",  X"08",  X"30",  X"08",  X"01",
  X"A0",  X"58",  X"FF",  X"1D",  X"00",  X"08",  X"00",  X"A0",
  X"00",  X"09",  X"00",  X"11",  X"0E",  X"00",  X"01",  X"18",
  X"0C",  X"00",  X"4D",  X"00",  X"18",  X"18",  X"18",  X"0D",
  X"F4",  X"0A",  X"08",  X"01",  X"08",  X"00",  X"32",  X"84",
  X"00",  X"06",  X"32",  X"08",  X"84",  X"08",  X"01",  X"98",
  X"08",  X"84",  X"84",  X"08",  X"01",  X"A0",  X"00",  X"1A",
  X"00",  X"09",  X"10",  X"18",  X"18",  X"01",  X"10",  X"12",
  X"00",  X"10",  X"18",  X"18",  X"0A",  X"F6",  X"00",  X"0C",
  X"0D",  X"10",  X"18",  X"08",  X"18",  X"01",  X"10",  X"F3",
  X"10",  X"08",  X"1A",  X"30",  X"34",  X"04",  X"00",  X"04",
  X"FE",  X"FF",  X"00",  X"0A",  X"04",  X"00",  X"08",  X"00",
  X"00",  X"04",  X"FE",  X"0D",  X"00",  X"08",  X"00",  X"30",
  X"34",  X"00",  X"04",  X"07",  X"00",  X"00",  X"01",  X"FE",
  X"00",  X"00",  X"08",  X"00",  X"00",  X"01",  X"01",  X"30",
  X"3C",  X"14",  X"01",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"08",  X"10",  X"18",  X"20",  X"28",  X"30",  X"38",
  X"00",  X"17",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"01",  X"30",  X"3C",  X"15",  X"14",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"08",  X"10",  X"18",  X"20",
  X"28",  X"30",  X"38",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"27",  X"94",  X"00",  X"30",  X"74",  X"00",  X"20",  X"00",
  X"00",  X"00",  X"A0",  X"A0",  X"A0",  X"A0",  X"A0",  X"A0",
  X"A0",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"30",  X"74",  X"00",  X"68",  X"04",  X"64",  X"68",  X"A9",
  X"00",  X"30",  X"58",  X"00",  X"04",  X"10",  X"14",  X"18",
  X"1C",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"30",  X"3C",  X"00",  X"01",  X"FF",  X"03",  X"00",  X"00",
  X"00",  X"F9",  X"00",  X"30",  X"3C",  X"00",  X"FF",  X"03",
  X"00",  X"00",  X"01",  X"00",  X"F9",  X"00",  X"00",  X"30",
  X"58",  X"04",  X"00",  X"10",  X"14",  X"18",  X"1C",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"04",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"04",  X"02",  X"05",  X"00",  X"00",
  X"20",  X"1F",  X"03",  X"06",  X"00",  X"00",  X"14",  X"00",
  X"18",  X"04",  X"08",  X"00",  X"40",  X"00",  X"00",  X"00",
  X"00",  X"0F",  X"05",  X"08",  X"00",  X"40",  X"00",  X"00",
  X"00",  X"00",  X"06",  X"06",  X"03",  X"00",  X"A3",  X"00",
  X"00",  X"04",  X"03",  X"08",  X"02",  X"02",  X"08",  X"02",
  X"06",  X"08",  X"02",  X"04",  X"13",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"04",  X"14",  X"03",  X"00",  X"00",
  X"30",  X"1C",  X"00",  X"30",  X"18",  X"00",  X"15",  X"2D",
  X"00",  X"15",  X"13",  X"00",  X"00",  X"08",  X"10",  X"18",
  X"20",  X"28",  X"30",  X"38",  X"40",  X"48",  X"50",  X"58",
  X"60",  X"68",  X"70",  X"78",  X"80",  X"30",  X"18",  X"00",
  X"14",  X"13",  X"00",  X"00",  X"08",  X"10",  X"18",  X"20",
  X"28",  X"30",  X"38",  X"40",  X"48",  X"50",  X"58",  X"60",
  X"68",  X"70",  X"78",  X"80",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"08",  X"00",  X"08",  X"00",  X"08",  X"00",
  X"10",  X"00",  X"26",  X"94",  X"28",  X"5C",  X"00",  X"30",
  X"28",  X"00",  X"01",  X"00",  X"08",  X"00",  X"09",  X"30",
  X"20",  X"00",  X"08",  X"02",  X"00",  X"20",  X"00",  X"00",
  X"00",  X"17",  X"37",  X"F8",  X"00",  X"20",  X"00",  X"00",
  X"00",  X"30",  X"28",  X"00",  X"01",  X"00",  X"39",  X"00",
  X"A0",  X"31",  X"02",  X"50",  X"1F",  X"00",  X"17",  X"04",
  X"04",  X"31",  X"00",  X"D0",  X"0D",  X"0C",  X"02",  X"06",
  X"03",  X"0E",  X"0C",  X"0C",  X"0C",  X"0C",  X"00",  X"FC",
  X"01",  X"04",  X"0C",  X"0C",  X"00",  X"08",  X"01",  X"0C",
  X"08",  X"01",  X"02",  X"31",  X"50",  X"08",  X"0C",  X"08",
  X"08",  X"A0",  X"30",  X"2C",  X"04",  X"18",  X"40",  X"2C",
  X"00",  X"02",  X"01",  X"02",  X"31",  X"50",  X"11",  X"00",
  X"34",  X"32",  X"32",  X"32",  X"32",  X"D0",  X"54",  X"58",
  X"1D",  X"D4",  X"13",  X"01",  X"11",  X"00",  X"00",  X"06",
  X"08",  X"00",  X"00",  X"00",  X"08",  X"18",  X"00",  X"19",
  X"00",  X"00",  X"05",  X"11",  X"00",  X"00",  X"11",  X"FF",
  X"11",  X"0C",  X"00",  X"11",  X"00",  X"00",  X"00",  X"FB",
  X"0C",  X"00",  X"00",  X"DF",  X"11",  X"00",  X"DD",  X"13",
  X"0C",  X"00",  X"F4",  X"00",  X"08",  X"00",  X"C0",  X"C1",
  X"1F",  X"0F",  X"00",  X"18",  X"0F",  X"03",  X"0C",  X"30",
  X"34",  X"00",  X"70",  X"00",  X"30",  X"50",  X"00",  X"40",
  X"00",  X"39",  X"01",  X"06",  X"FC",  X"00",  X"08",  X"33",
  X"00",  X"10",  X"00",  X"08",  X"FC",  X"08",  X"02",  X"01",
  X"0C",  X"05",  X"00",  X"08",  X"26",  X"00",  X"15",  X"01",
  X"30",  X"34",  X"00",  X"02",  X"01",  X"11",  X"F8",  X"00",
  X"08",  X"19",  X"00",  X"08",  X"01",  X"10",  X"30",  X"50",
  X"00",  X"02",  X"01",  X"0D",  X"EA",  X"00",  X"08",  X"0B",
  X"00",  X"FA",  X"01",  X"30",  X"2C",  X"00",  X"10",  X"10",
  X"0F",  X"04",  X"06",  X"08",  X"00",  X"30",  X"48",  X"01",
  X"00",  X"08",  X"00",  X"A0",  X"32",  X"60",  X"18",  X"00",
  X"06",  X"00",  X"02",  X"00",  X"19",  X"08",  X"08",  X"00",
  X"A0",  X"32",  X"64",  X"00",  X"05",  X"00",  X"00",  X"18",
  X"08",  X"08",  X"02",  X"A0",  X"32",  X"6C",  X"00",  X"05",
  X"00",  X"00",  X"18",  X"08",  X"08",  X"02",  X"A0",  X"32",
  X"68",  X"00",  X"05",  X"00",  X"00",  X"18",  X"08",  X"08",
  X"02",  X"A0",  X"32",  X"70",  X"00",  X"05",  X"00",  X"00",
  X"18",  X"08",  X"08",  X"02",  X"A0",  X"32",  X"74",  X"00",
  X"05",  X"00",  X"00",  X"18",  X"08",  X"08",  X"02",  X"A0",
  X"32",  X"78",  X"00",  X"05",  X"00",  X"00",  X"18",  X"08",
  X"08",  X"02",  X"A0",  X"32",  X"7C",  X"18",  X"00",  X"06",
  X"00",  X"02",  X"00",  X"19",  X"08",  X"08",  X"00",  X"00",
  X"27",  X"6C",  X"00",  X"00",  X"00",  X"00",  X"00",  X"27",
  X"F0",  X"00",  X"00",  X"27",  X"5C",  X"00",  X"00",  X"00",
  X"18",  X"03",  X"03",  X"07",  X"00",  X"00",  X"1C",  X"00",
  X"06",  X"00",  X"37",  X"00",  X"E2",  X"00",  X"40",  X"79",
  X"00",  X"01",  X"00",  X"00",  X"04",  X"14",  X"03",  X"14",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"04",  X"08",
  X"00",  X"08",  X"00",  X"00",  X"18",  X"03",  X"03",  X"08",
  X"00",  X"30",  X"44",  X"03",  X"00",  X"00",  X"08",  X"30",
  X"44",  X"02",  X"00",  X"00",  X"24",  X"14",  X"1F",  X"30",
  X"3C",  X"00",  X"01",  X"30",  X"38",  X"00",  X"30",  X"40",
  X"02",  X"00",  X"08",  X"00",  X"08",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"18",  X"03",  X"03",
  X"06",  X"00",  X"00",  X"08",  X"02",  X"00",  X"00",  X"27",
  X"A0",  X"00",  X"A0",  X"2C",  X"2C",  X"C0",  X"C0",  X"11",
  X"0B",  X"00",  X"00",  X"00",  X"04",  X"04",  X"00",  X"00",
  X"11",  X"FA",  X"00",  X"08",  X"00",  X"40",  X"60",  X"64",
  X"68",  X"74",  X"78",  X"80",  X"88",  X"00",  X"6C",  X"90",
  X"98",  X"A0",  X"A8",  X"30",  X"1C",  X"3C",  X"B0",  X"1C",
  X"01",  X"10",  X"13",  X"13",  X"00",  X"01",  X"30",  X"3C",
  X"03",  X"02",  X"FF",  X"00",  X"00",  X"00",  X"08",  X"10",
  X"18",  X"20",  X"28",  X"30",  X"38",  X"00",  X"08",  X"15",
  X"32",  X"5C",  X"00",  X"00",  X"04",  X"00",  X"00",  X"F8",
  X"3C",  X"30",  X"1C",  X"00",  X"02",  X"10",  X"30",  X"38",
  X"02",  X"02",  X"00",  X"01",  X"20",  X"01",  X"30",  X"3C",
  X"03",  X"02",  X"FF",  X"00",  X"6C",  X"00",  X"90",  X"98",
  X"A0",  X"A8",  X"74",  X"78",  X"80",  X"88",  X"60",  X"64",
  X"68",  X"00",  X"00",  X"08",  X"10",  X"18",  X"20",  X"28",
  X"30",  X"38",  X"0F",  X"00",  X"6C",  X"00",  X"90",  X"98",
  X"A0",  X"A8",  X"74",  X"78",  X"80",  X"88",  X"60",  X"64",
  X"68",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"40",
  X"38",  X"04",  X"14",  X"74",  X"78",  X"80",  X"88",  X"00",
  X"6C",  X"30",  X"1C",  X"3C",  X"B0",  X"1C",  X"80",  X"01",
  X"10",  X"13",  X"13",  X"00",  X"01",  X"30",  X"3C",  X"03",
  X"02",  X"FF",  X"00",  X"00",  X"00",  X"08",  X"10",  X"18",
  X"20",  X"28",  X"30",  X"38",  X"00",  X"08",  X"15",  X"32",
  X"5C",  X"00",  X"00",  X"04",  X"00",  X"00",  X"F8",  X"3C",
  X"30",  X"1C",  X"30",  X"18",  X"03",  X"08",  X"00",  X"38",
  X"04",  X"03",  X"03",  X"02",  X"06",  X"B0",  X"03",  X"03",
  X"30",  X"18",  X"00",  X"02",  X"10",  X"30",  X"38",  X"02",
  X"02",  X"00",  X"01",  X"19",  X"01",  X"30",  X"3C",  X"03",
  X"02",  X"FF",  X"00",  X"6C",  X"00",  X"74",  X"78",  X"80",
  X"88",  X"00",  X"00",  X"08",  X"10",  X"18",  X"20",  X"28",
  X"30",  X"38",  X"08",  X"00",  X"6C",  X"00",  X"74",  X"78",
  X"80",  X"88",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"08",  X"00",  X"00",  X"05",  X"08",  X"08",  X"18",  X"01",
  X"08",  X"01",  X"0C",  X"FF",  X"09",  X"07",  X"0C",  X"01",
  X"07",  X"F3",  X"05",  X"00",  X"08",  X"0A",  X"08",  X"00",
  X"03",  X"08",  X"08",  X"18",  X"09",  X"08",  X"01",  X"0C",
  X"FF",  X"0A",  X"07",  X"0D",  X"01",  X"0F",  X"F3",  X"03",
  X"00",  X"08",  X"0B",  X"04",  X"00",  X"0B",  X"0B",  X"0C",
  X"08",  X"3F",  X"F0",  X"08",  X"04",  X"0B",  X"0A",  X"08",
  X"09",  X"2D",  X"08",  X"F0",  X"A0",  X"2C",  X"A8",  X"FC",
  X"FF",  X"08",  X"FC",  X"00",  X"FC",  X"00",  X"FF",  X"FC",
  X"00",  X"08",  X"00",  X"A0",  X"08",  X"00",  X"00",  X"00",
  X"10",  X"00",  X"00",  X"01",  X"00",  X"10",  X"18",  X"1C",
  X"08",  X"00",  X"18",  X"00",  X"52",  X"0F",  X"00",  X"0C",
  X"00",  X"18",  X"20",  X"F4",  X"7C",  X"1E",  X"0F",  X"00",
  X"18",  X"3C",  X"54",  X"20",  X"1E",  X"0F",  X"00",  X"18",
  X"58",  X"58",  X"14",  X"1E",  X"0F",  X"00",  X"18",  X"74",
  X"50",  X"60",  X"1E",  X"0F",  X"00",  X"18",  X"90",  X"94",
  X"60",  X"1E",  X"0F",  X"00",  X"18",  X"AC",  X"D8",  X"C0",
  X"1E",  X"0F",  X"00",  X"18",  X"C8",  X"7C",  X"54",  X"1E",
  X"0F",  X"00",  X"18",  X"E4",  X"B4",  X"AC",  X"1E",  X"0F",
  X"00",  X"18",  X"00",  X"44",  X"44",  X"1E",  X"0F",  X"00",
  X"18",  X"1C",  X"6C",  X"48",  X"1E",  X"0F",  X"00",  X"18",
  X"38",  X"98",  X"34",  X"1E",  X"0F",  X"00",  X"10",  X"7C",
  X"B0",  X"20",  X"00",  X"18",  X"90",  X"BC",  X"50",  X"1E",
  X"0F",  X"00",  X"18",  X"AC",  X"F0",  X"54",  X"1E",  X"0F",
  X"00",  X"18",  X"C8",  X"28",  X"2C",  X"1E",  X"0F",  X"00",
  X"10",  X"E4",  X"38",  X"1C",  X"00",  X"10",  X"F8",  X"40",
  X"1C",  X"00",  X"18",  X"0C",  X"48",  X"D8",  X"1E",  X"0F",
  X"00",  X"10",  X"28",  X"04",  X"18",  X"00",  X"10",  X"3C",
  X"08",  X"18",  X"00",  X"18",  X"50",  X"0C",  X"40",  X"1E",
  X"0F",  X"00",  X"18",  X"6C",  X"94",  X"38",  X"1E",  X"0F",
  X"00",  X"14",  X"88",  X"B0",  X"54",  X"1E",  X"1F",  X"10",
  X"A0",  X"EC",  X"2C",  X"00",  X"18",  X"B4",  X"04",  X"60",
  X"1E",  X"0F",  X"00",  X"10",  X"D0",  X"48",  X"2C",  X"00",
  X"18",  X"E4",  X"60",  X"38",  X"1E",  X"0F",  X"00",  X"10",
  X"00",  X"7C",  X"34",  X"00",  X"18",  X"14",  X"9C",  X"F4",
  X"1E",  X"0F",  X"00",  X"18",  X"30",  X"74",  X"34",  X"1E",
  X"0F",  X"00",  X"18",  X"4C",  X"8C",  X"18",  X"1E",  X"0F",
  X"00",  X"18",  X"68",  X"88",  X"04",  X"1E",  X"0F",  X"00",
  X"18",  X"84",  X"70",  X"5C",  X"1E",  X"0F",  X"00",  X"10",
  X"A0",  X"B0",  X"18",  X"00",  X"10",  X"B4",  X"B4",  X"18",
  X"00",  X"18",  X"C8",  X"B8",  X"24",  X"1E",  X"0F",  X"00",
  X"10",  X"E4",  X"C0",  X"18",  X"00",  X"18",  X"F8",  X"C4",
  X"24",  X"1E",  X"0F",  X"00",  X"18",  X"14",  X"CC",  X"24",
  X"1E",  X"0F",  X"00",  X"10",  X"30",  X"D4",  X"18",  X"00",
  X"14",  X"44",  X"D8",  X"20",  X"1E",  X"1F",  X"18",  X"5C",
  X"E0",  X"8C",  X"1E",  X"0F",  X"00",  X"18",  X"78",  X"50",
  X"6C",  X"1E",  X"0F",  X"00",  X"18",  X"94",  X"A0",  X"50",
  X"1E",  X"0F",  X"00",  X"14",  X"B0",  X"D4",  X"1C",  X"1E",
  X"1F",  X"14",  X"C8",  X"D8",  X"EC",  X"1E",  X"1F",  X"18",
  X"E0",  X"AC",  X"9C",  X"1E",  X"0F",  X"00",  X"18",  X"FC",
  X"2C",  X"20",  X"1E",  X"0F",  X"00",  X"14",  X"18",  X"30",
  X"E4",  X"1E",  X"1F",  X"14",  X"30",  X"FC",  X"E0",  X"1E",
  X"1F",  X"10",  X"48",  X"C4",  X"0C",  X"00",  X"10",  X"5C",
  X"BC",  X"0C",  X"00",  X"10",  X"70",  X"B4",  X"0C",  X"00",
  X"18",  X"84",  X"AC",  X"68",  X"1E",  X"0F",  X"00",  X"10",
  X"A0",  X"F8",  X"24",  X"00",  X"18",  X"B4",  X"08",  X"60",
  X"1E",  X"0F",  X"00",  X"18",  X"D0",  X"4C",  X"F0",  X"1E",
  X"0F",  X"00",  X"18",  X"EC",  X"20",  X"FC",  X"1E",  X"0F",
  X"00",  X"18",  X"08",  X"00",  X"50",  X"1E",  X"0F",  X"00",
  X"18",  X"24",  X"34",  X"DC",  X"1E",  X"0F",  X"00",  X"10",
  X"40",  X"F4",  X"2C",  X"00",  X"10",  X"54",  X"0C",  X"84",
  X"00",  X"10",  X"68",  X"7C",  X"E4",  X"00",  X"18",  X"7C",
  X"4C",  X"74",  X"1E",  X"0F",  X"00",  X"10",  X"98",  X"A4",
  X"9C",  X"68",  X"18",  X"AC",  X"2C",  X"10",  X"1E",  X"0F",
  X"00",  X"18",  X"C8",  X"20",  X"AC",  X"1E",  X"0F",  X"00",
  X"10",  X"E4",  X"B0",  X"40",  X"00",  X"18",  X"F8",  X"DC",
  X"A8",  X"1E",  X"0F",  X"00",  X"18",  X"14",  X"68",  X"30",
  X"1E",  X"0F",  X"00",  X"18",  X"30",  X"7C",  X"B4",  X"1E",
  X"0F",  X"00",  X"18",  X"4C",  X"14",  X"34",  X"1E",  X"0F",
  X"00",  X"18",  X"68",  X"2C",  X"20",  X"1E",  X"0F",  X"00",
  X"18",  X"84",  X"30",  X"24",  X"1E",  X"0F",  X"00",  X"18",
  X"A0",  X"38",  X"E8",  X"1E",  X"0F",  X"00",  X"18",  X"BC",
  X"04",  X"14",  X"1E",  X"0F",  X"00",  X"18",  X"D8",  X"FC",
  X"D0",  X"1E",  X"0F",  X"00",  X"18",  X"F4",  X"B0",  X"F8",
  X"1E",  X"0F",  X"00",  X"18",  X"10",  X"8C",  X"8C",  X"1E",
  X"0F",  X"00",  X"18",  X"2C",  X"FC",  X"28",  X"1E",  X"0F",
  X"00",  X"18",  X"48",  X"08",  X"04",  X"1E",  X"0F",  X"00",
  X"10",  X"64",  X"F0",  X"34",  X"00",  X"10",  X"78",  X"10",
  X"28",  X"00",  X"10",  X"8C",  X"24",  X"1C",  X"00",  X"18",
  X"A0",  X"2C",  X"58",  X"1E",  X"0F",  X"00",  X"18",  X"BC",
  X"68",  X"58",  X"1E",  X"0F",  X"00",  X"18",  X"D8",  X"A4",
  X"50",  X"1E",  X"0F",  X"00",  X"10",  X"F4",  X"D8",  X"E8",
  X"00",  X"18",  X"08",  X"AC",  X"94",  X"1E",  X"0F",  X"00",
  X"18",  X"24",  X"24",  X"48",  X"1E",  X"0F",  X"00",  X"18",
  X"40",  X"50",  X"A0",  X"1E",  X"0F",  X"00",  X"18",  X"5C",
  X"D4",  X"40",  X"1E",  X"0F",  X"00",  X"18",  X"78",  X"F8",
  X"70",  X"1E",  X"0F",  X"00",  X"10",  X"94",  X"4C",  X"1C",
  X"00",  X"18",  X"A8",  X"54",  X"44",  X"1E",  X"0F",  X"00",
  X"18",  X"C4",  X"7C",  X"48",  X"1E",  X"0F",  X"00",  X"18",
  X"E0",  X"A8",  X"48",  X"1E",  X"0F",  X"00",  X"10",  X"FC",
  X"1C",  X"08",  X"00",  X"10",  X"10",  X"10",  X"14",  X"00",
  X"10",  X"24",  X"10",  X"08",  X"00",  X"14",  X"38",  X"04",
  X"1C",  X"1E",  X"1F",  X"18",  X"50",  X"08",  X"5C",  X"1E",
  X"0F",  X"00",  X"10",  X"6C",  X"48",  X"3C",  X"00",  X"18",
  X"80",  X"70",  X"78",  X"1E",  X"0F",  X"00",  X"10",  X"9C",
  X"CC",  X"50",  X"00",  X"10",  X"B0",  X"08",  X"34",  X"00",
  X"18",  X"C4",  X"F8",  X"88",  X"1E",  X"0F",  X"00",  X"10",
  X"E0",  X"64",  X"1C",  X"00",  X"18",  X"F4",  X"6C",  X"20",
  X"1E",  X"0F",  X"00",  X"10",  X"10",  X"A8",  X"10",  X"00",
  X"18",  X"24",  X"A4",  X"34",  X"1E",  X"0F",  X"00",  X"18",
  X"40",  X"BC",  X"2C",  X"1E",  X"0F",  X"00",  X"18",  X"5C",
  X"CC",  X"2C",  X"1E",  X"0F",  X"00",  X"18",  X"78",  X"DC",
  X"2C",  X"1E",  X"0F",  X"00",  X"18",  X"94",  X"EC",  X"2C",
  X"1E",  X"0F",  X"00",  X"18",  X"B0",  X"FC",  X"2C",  X"1E",
  X"0F",  X"00",  X"18",  X"CC",  X"0C",  X"2C",  X"1E",  X"0F",
  X"00",  X"18",  X"E8",  X"1C",  X"34",  X"1E",  X"0F",  X"00",
  X"18",  X"04",  X"E0",  X"4C",  X"1E",  X"0F",  X"00",  X"10",
  X"20",  X"80",  X"0C",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"02",  X"FF",  X"00",  X"00",  X"02",  X"FF",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"02",  X"00",  X"01",  X"02",  X"03",
  X"04",  X"06",  X"01",  X"02",  X"04",  X"08",  X"10",  X"20",
  X"40",  X"80",  X"00",  X"00",  X"00",  X"00",  X"01",  X"02",
  X"04",  X"08",  X"10",  X"20",  X"40",  X"80",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"01",  X"02",  X"04",
  X"08",  X"10",  X"20",  X"00",  X"00",  X"00",  X"02",  X"00",
  X"01",  X"02",  X"03",  X"04",  X"06",  X"01",  X"02",  X"04",
  X"08",  X"10",  X"20",  X"00",  X"20",  X"00",  X"34",  X"00",
  X"01",  X"02",  X"04",  X"08",  X"10",  X"20",  X"40",  X"80",
  X"00",  X"00",  X"00",  X"00",  X"01",  X"02",  X"04",  X"08",
  X"10",  X"20",  X"40",  X"80",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"02",
  X"00",  X"01",  X"02",  X"03",  X"04",  X"06",  X"01",  X"02",
  X"04",  X"08",  X"10",  X"20",  X"40",  X"80",  X"00",  X"00",
  X"00",  X"00",  X"01",  X"02",  X"04",  X"08",  X"10",  X"20",
  X"40",  X"80",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"01",  X"02",  X"04",  X"08",  X"10",  X"20",  X"40",
  X"80",  X"00",  X"00",  X"00",  X"00",  X"01",  X"02",  X"04",
  X"08",  X"10",  X"20",  X"40",  X"80",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"02",
  X"00",  X"01",  X"02",  X"03",  X"04",  X"06",  X"01",  X"02",
  X"04",  X"08",  X"10",  X"20",  X"B8",  X"1F",  X"00",  X"00",
  X"00",  X"02",  X"00",  X"01",  X"02",  X"03",  X"04",  X"06",
  X"01",  X"02",  X"04",  X"08",  X"10",  X"20",  X"01",  X"02",
  X"04",  X"08",  X"10",  X"20",  X"40",  X"80",  X"00",  X"00",
  X"00",  X"00",  X"01",  X"02",  X"04",  X"08",  X"10",  X"20",
  X"40",  X"80",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"F8",  X"00",  X"00",  X"00",  X"33",  X"37",
  X"42",  X"46",  X"00",  X"00",  X"00",  X"00",  X"33",  X"37",
  X"62",  X"66",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"6C",  X"00",  X"00",  X"00",  X"30",  X"30",
  X"30",  X"30",  X"20",  X"20",  X"20",  X"20",  X"54",  X"00",
  X"4A",  X"00",  X"55",  X"00",  X"49",  X"00",  X"69",  X"79",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"A7",  X"61",
  X"28",  X"B3",  X"13",  X"FB",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"2D",  X"39",
  X"00",  X"00",  X"80",  X"48",  X"48",  X"48",  X"48",  X"48",
  X"48",  X"48",  X"48",  X"48",  X"7F",  X"7F",  X"38",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"80",  X"00",  X"D0",  X"00",
  X"84",  X"00",  X"65",  X"00",  X"5F",  X"00",  X"76",  X"00",
  X"94",  X"00",  X"9C",  X"00",  X"C4",  X"00",  X"F5",  X"00",
  X"79",  X"00",  X"57",  X"00",  X"6D",  X"00",  X"E4",  X"00",
  X"1D",  X"40",  X"E4",  X"50",  X"CF",  X"92",  X"02",  X"F6",
  X"43",  X"B4",  X"79",  X"00",  X"B5",  X"17",  X"03",  X"F5",
  X"48",  X"32",  X"DD",  X"3C",  X"B2",  X"BC",  X"23",  X"33",
  X"FD",  X"3D",  X"08",  X"9D",  X"28",  X"43",  X"05",  X"19",
  X"7D",  X"00",  X"A0",  X"9F",  X"00",  X"57",  X"00",  X"08",
  X"00",  X"A0",  X"6D",  X"00",  X"08",  X"00",  X"00",  X"00",
  X"01",  X"00",  X"00",  X"00",  X"F8",  X"00",  X"00",  X"E4",
  X"B0",  X"7C",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"30",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"01",  X"CD",  X"6D",  X"05",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"48",  X"48",  X"50",  X"50",
  X"58",  X"58",  X"60",  X"60",  X"68",  X"68",  X"70",  X"70",
  X"78",  X"78",  X"80",  X"80",  X"88",  X"88",  X"90",  X"90",
  X"98",  X"98",  X"A0",  X"A0",  X"A8",  X"A8",  X"B0",  X"B0",
  X"B8",  X"B8",  X"C0",  X"C0",  X"C8",  X"C8",  X"D0",  X"D0",
  X"D8",  X"D8",  X"E0",  X"E0",  X"E8",  X"E8",  X"F0",  X"F0",
  X"F8",  X"F8",  X"00",  X"00",  X"08",  X"08",  X"10",  X"10",
  X"18",  X"18",  X"20",  X"20",  X"28",  X"28",  X"30",  X"30",
  X"38",  X"38",  X"40",  X"40",  X"48",  X"48",  X"50",  X"50",
  X"58",  X"58",  X"60",  X"60",  X"68",  X"68",  X"70",  X"70",
  X"78",  X"78",  X"80",  X"80",  X"88",  X"88",  X"90",  X"90",
  X"98",  X"98",  X"A0",  X"A0",  X"A8",  X"A8",  X"B0",  X"B0",
  X"B8",  X"B8",  X"C0",  X"C0",  X"C8",  X"C8",  X"D0",  X"D0",
  X"D8",  X"D8",  X"E0",  X"E0",  X"E8",  X"E8",  X"F0",  X"F0",
  X"F8",  X"F8",  X"00",  X"00",  X"08",  X"08",  X"10",  X"10",
  X"18",  X"18",  X"20",  X"20",  X"28",  X"28",  X"30",  X"30",
  X"38",  X"38",  X"40",  X"40",  X"48",  X"48",  X"50",  X"50",
  X"58",  X"58",  X"60",  X"60",  X"68",  X"68",  X"70",  X"70",
  X"78",  X"78",  X"80",  X"80",  X"88",  X"88",  X"90",  X"90",
  X"98",  X"98",  X"A0",  X"A0",  X"A8",  X"A8",  X"B0",  X"B0",
  X"B8",  X"B8",  X"C0",  X"C0",  X"C8",  X"C8",  X"D0",  X"D0",
  X"D8",  X"D8",  X"E0",  X"E0",  X"E8",  X"E8",  X"F0",  X"F0",
  X"F8",  X"F8",  X"00",  X"00",  X"08",  X"08",  X"10",  X"10",
  X"18",  X"18",  X"20",  X"20",  X"28",  X"28",  X"30",  X"30",
  X"38",  X"38",  X"40",  X"40",  X"48",  X"48",  X"50",  X"50",
  X"58",  X"58",  X"60",  X"60",  X"68",  X"68",  X"70",  X"70",
  X"78",  X"78",  X"80",  X"80",  X"88",  X"88",  X"90",  X"90",
  X"98",  X"98",  X"A0",  X"A0",  X"A8",  X"A8",  X"B0",  X"B0",
  X"B8",  X"B8",  X"C0",  X"C0",  X"C8",  X"C8",  X"D0",  X"D0",
  X"D8",  X"D8",  X"E0",  X"E0",  X"E8",  X"E8",  X"F0",  X"F0",
  X"F8",  X"F8",  X"00",  X"00",  X"08",  X"08",  X"10",  X"10",
  X"18",  X"18",  X"20",  X"20",  X"28",  X"28",  X"30",  X"30",
  X"38",  X"38",  X"40",  X"40",  X"00",  X"FF",  X"00",  X"58",
  X"00",  X"00",  X"00",  X"02",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"CC",  X"00",  X"00",  X"00",
  X"02",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"01",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"78",  X"78",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"08",  X"07",
  X"06",  X"03",  X"00",  X"D0",  X"10",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  others => X"00" );


constant ram01 : ram_type := (
  X"00",  X"00",  X"23",  X"00",  X"00",  X"00",  X"27",  X"20",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"23",  X"00",  X"00",  X"00",  X"20",  X"00",
  X"00",  X"00",  X"20",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"00",  X"00",  X"27",  X"20",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"25",  X"00",
  X"20",  X"00",  X"25",  X"00",  X"20",  X"00",  X"25",  X"00",
  X"20",  X"00",  X"25",  X"00",  X"20",  X"00",  X"25",  X"00",
  X"20",  X"00",  X"25",  X"00",  X"20",  X"00",  X"25",  X"00",
  X"20",  X"00",  X"25",  X"00",  X"20",  X"00",  X"25",  X"00",
  X"20",  X"00",  X"25",  X"00",  X"20",  X"00",  X"25",  X"00",
  X"20",  X"00",  X"25",  X"00",  X"20",  X"00",  X"25",  X"00",
  X"20",  X"00",  X"25",  X"00",  X"20",  X"00",  X"25",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"22",  X"00",  X"00",  X"23",  X"00",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"00",  X"00",  X"22",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"BF",  X"00",  X"A2",  X"00",  X"E1",  X"00",  X"C0",  X"E0",
  X"FF",  X"80",  X"00",  X"21",  X"00",  X"22",  X"00",  X"22",
  X"00",  X"23",  X"00",  X"00",  X"22",  X"01",  X"00",  X"29",
  X"00",  X"01",  X"00",  X"22",  X"00",  X"E0",  X"00",  X"BF",
  X"00",  X"22",  X"60",  X"00",  X"00",  X"62",  X"00",  X"00",
  X"E0",  X"A0",  X"80",  X"A0",  X"BF",  X"40",  X"00",  X"00",
  X"62",  X"60",  X"60",  X"40",  X"C0",  X"40",  X"00",  X"40",
  X"40",  X"FF",  X"60",  X"00",  X"60",  X"60",  X"00",  X"20",
  X"00",  X"FB",  X"20",  X"20",  X"22",  X"E0",  X"00",  X"BF",
  X"E0",  X"00",  X"BF",  X"00",  X"60",  X"60",  X"00",  X"00",
  X"00",  X"00",  X"20",  X"FB",  X"62",  X"00",  X"21",  X"60",
  X"00",  X"21",  X"00",  X"60",  X"60",  X"00",  X"00",  X"40",
  X"00",  X"E0",  X"00",  X"BF",  X"E0",  X"00",  X"E0",  X"00",
  X"BF",  X"A0",  X"A0",  X"A0",  X"A0",  X"A0",  X"A0",  X"BF",
  X"A0",  X"BF",  X"BF",  X"00",  X"A2",  X"A0",  X"00",  X"01",
  X"00",  X"00",  X"BF",  X"00",  X"63",  X"00",  X"62",  X"BF",
  X"00",  X"00",  X"BF",  X"00",  X"00",  X"E0",  X"00",  X"BF",
  X"00",  X"63",  X"00",  X"00",  X"00",  X"E0",  X"00",  X"BF",
  X"A0",  X"A0",  X"62",  X"60",  X"00",  X"00",  X"A0",  X"40",
  X"A0",  X"80",  X"A0",  X"FF",  X"A3",  X"C0",  X"60",  X"00",
  X"00",  X"A0",  X"40",  X"A0",  X"A2",  X"A0",  X"A2",  X"00",
  X"C0",  X"80",  X"A0",  X"A0",  X"40",  X"A0",  X"62",  X"7F",
  X"A0",  X"62",  X"A0",  X"62",  X"60",  X"00",  X"3F",  X"60",
  X"60",  X"00",  X"00",  X"A0",  X"40",  X"A0",  X"80",  X"A0",
  X"FF",  X"A3",  X"C0",  X"60",  X"00",  X"00",  X"A0",  X"40",
  X"60",  X"62",  X"60",  X"00",  X"3F",  X"60",  X"60",  X"FF",
  X"00",  X"00",  X"E0",  X"00",  X"BF",  X"A0",  X"A0",  X"A0",
  X"A0",  X"BF",  X"A0",  X"62",  X"A0",  X"80",  X"A0",  X"62",
  X"A0",  X"62",  X"61",  X"00",  X"00",  X"A0",  X"21",  X"62",
  X"BF",  X"00",  X"00",  X"A0",  X"62",  X"A0",  X"62",  X"7F",
  X"BF",  X"A0",  X"00",  X"C0",  X"40",  X"40",  X"80",  X"A0",
  X"62",  X"60",  X"A0",  X"62",  X"A0",  X"62",  X"A0",  X"62",
  X"80",  X"3F",  X"60",  X"60",  X"00",  X"00",  X"A0",  X"61",
  X"A0",  X"62",  X"BF",  X"60",  X"BF",  X"20",  X"BF",  X"A0",
  X"C0",  X"00",  X"00",  X"20",  X"60",  X"60",  X"FF",  X"00",
  X"A0",  X"62",  X"60",  X"00",  X"00",  X"A0",  X"40",  X"A0",
  X"80",  X"A0",  X"00",  X"00",  X"C0",  X"60",  X"A0",  X"FF",
  X"00",  X"00",  X"E0",  X"00",  X"BF",  X"A0",  X"A0",  X"00",
  X"A1",  X"40",  X"A0",  X"40",  X"20",  X"60",  X"A0",  X"61",
  X"A0",  X"62",  X"A0",  X"62",  X"A0",  X"40",  X"00",  X"A0",
  X"60",  X"00",  X"E0",  X"00",  X"BF",  X"A0",  X"A0",  X"00",
  X"A3",  X"40",  X"A0",  X"40",  X"20",  X"60",  X"A0",  X"40",
  X"20",  X"40",  X"BF",  X"00",  X"00",  X"A0",  X"40",  X"BF",
  X"60",  X"80",  X"60",  X"BF",  X"60",  X"BF",  X"20",  X"BF",
  X"A0",  X"00",  X"00",  X"20",  X"60",  X"60",  X"FF",  X"00",
  X"A0",  X"40",  X"03",  X"A2",  X"60",  X"A0",  X"40",  X"20",
  X"60",  X"00",  X"E0",  X"00",  X"BF",  X"00",  X"63",  X"40",
  X"60",  X"00",  X"63",  X"40",  X"00",  X"63",  X"40",  X"00",
  X"A1",  X"00",  X"A1",  X"00",  X"FE",  X"00",  X"00",  X"E0",
  X"00",  X"BF",  X"A0",  X"A0",  X"00",  X"A2",  X"40",  X"A0",
  X"40",  X"40",  X"A0",  X"40",  X"60",  X"A0",  X"40",  X"3F",
  X"60",  X"00",  X"61",  X"20",  X"20",  X"00",  X"00",  X"62",
  X"20",  X"20",  X"00",  X"A0",  X"40",  X"A0",  X"80",  X"A0",
  X"A0",  X"60",  X"A0",  X"40",  X"A0",  X"80",  X"A0",  X"A0",
  X"60",  X"00",  X"E0",  X"00",  X"BF",  X"A0",  X"A0",  X"A0",
  X"40",  X"A0",  X"80",  X"A0",  X"20",  X"A0",  X"00",  X"00",
  X"C0",  X"60",  X"00",  X"E0",  X"00",  X"BF",  X"A0",  X"00",
  X"63",  X"FF",  X"00",  X"A0",  X"60",  X"00",  X"FF",  X"00",
  X"A0",  X"00",  X"FF",  X"00",  X"00",  X"E0",  X"00",  X"BF",
  X"00",  X"63",  X"FF",  X"00",  X"00",  X"63",  X"40",  X"BF",
  X"20",  X"BF",  X"00",  X"00",  X"00",  X"20",  X"20",  X"20",
  X"C0",  X"00",  X"40",  X"00",  X"BE",  X"22",  X"BF",  X"FF",
  X"63",  X"BF",  X"BF",  X"3F",  X"BF",  X"BF",  X"00",  X"BF",
  X"00",  X"00",  X"02",  X"BF",  X"BF",  X"40",  X"E0",  X"00",
  X"BE",  X"00",  X"62",  X"22",  X"BF",  X"FF",  X"63",  X"BF",
  X"BF",  X"3F",  X"BF",  X"BF",  X"BF",  X"00",  X"00",  X"02",
  X"BF",  X"BF",  X"40",  X"E0",  X"00",  X"BF",  X"00",  X"21",
  X"21",  X"00",  X"60",  X"61",  X"20",  X"00",  X"61",  X"20",
  X"60",  X"00",  X"00",  X"20",  X"00",  X"60",  X"20",  X"60",
  X"A0",  X"60",  X"E0",  X"21",  X"00",  X"00",  X"20",  X"C0",
  X"40",  X"21",  X"20",  X"00",  X"00",  X"60",  X"A0",  X"60",
  X"20",  X"00",  X"20",  X"20",  X"21",  X"E0",  X"00",  X"00",
  X"21",  X"20",  X"00",  X"21",  X"61",  X"00",  X"61",  X"20",
  X"21",  X"21",  X"FF",  X"20",  X"21",  X"40",  X"00",  X"60",
  X"A0",  X"21",  X"60",  X"00",  X"20",  X"20",  X"20",  X"21",
  X"E0",  X"00",  X"FF",  X"61",  X"20",  X"3F",  X"E0",  X"00",
  X"00",  X"00",  X"62",  X"C0",  X"12",  X"40",  X"00",  X"00",
  X"00",  X"62",  X"C0",  X"00",  X"40",  X"00",  X"BF",  X"20",
  X"60",  X"60",  X"00",  X"20",  X"7F",  X"20",  X"00",  X"00",
  X"A0",  X"00",  X"00",  X"01",  X"00",  X"21",  X"00",  X"20",
  X"00",  X"60",  X"40",  X"60",  X"80",  X"01",  X"20",  X"A0",
  X"A0",  X"A0",  X"FF",  X"80",  X"E0",  X"20",  X"A0",  X"E0",
  X"60",  X"00",  X"01",  X"A0",  X"E0",  X"00",  X"60",  X"E0",
  X"3F",  X"00",  X"60",  X"00",  X"00",  X"00",  X"00",  X"62",
  X"E0",  X"60",  X"7F",  X"00",  X"40",  X"6F",  X"70",  X"00",
  X"01",  X"00",  X"3F",  X"00",  X"00",  X"C0",  X"80",  X"00",
  X"00",  X"40",  X"00",  X"A2",  X"60",  X"60",  X"BF",  X"80",
  X"60",  X"01",  X"00",  X"01",  X"00",  X"E0",  X"20",  X"20",
  X"60",  X"00",  X"20",  X"60",  X"00",  X"20",  X"60",  X"60",
  X"00",  X"20",  X"60",  X"01",  X"61",  X"20",  X"20",  X"20",
  X"00",  X"60",  X"40",  X"E0",  X"C0",  X"00",  X"A0",  X"00",
  X"20",  X"00",  X"A0",  X"A0",  X"C0",  X"00",  X"20",  X"A0",
  X"BF",  X"80",  X"60",  X"FF",  X"60",  X"3F",  X"20",  X"00",
  X"E0",  X"E0",  X"C0",  X"00",  X"60",  X"A0",  X"BF",  X"80",
  X"60",  X"00",  X"60",  X"E0",  X"00",  X"E0",  X"A1",  X"00",
  X"A0",  X"A0",  X"60",  X"00",  X"60",  X"A0",  X"20",  X"20",
  X"40",  X"60",  X"40",  X"00",  X"60",  X"00",  X"60",  X"40",
  X"00",  X"60",  X"60",  X"3F",  X"80",  X"FF",  X"60",  X"60",
  X"A0",  X"A0",  X"60",  X"A0",  X"60",  X"20",  X"20",  X"00",
  X"40",  X"FF",  X"60",  X"40",  X"00",  X"3F",  X"20",  X"00",
  X"40",  X"00",  X"60",  X"40",  X"00",  X"A0",  X"00",  X"E0",
  X"00",  X"A0",  X"A0",  X"40",  X"00",  X"E0",  X"A0",  X"BF",
  X"80",  X"60",  X"FF",  X"60",  X"A0",  X"A0",  X"80",  X"20",
  X"60",  X"20",  X"E0",  X"E0",  X"A0",  X"80",  X"A0",  X"00",
  X"A0",  X"A0",  X"80",  X"A0",  X"20",  X"E0",  X"A0",  X"60",
  X"00",  X"00",  X"A0",  X"E0",  X"00",  X"80",  X"A0",  X"60",
  X"A0",  X"00",  X"00",  X"A0",  X"E0",  X"00",  X"20",  X"FF",
  X"20",  X"A0",  X"40",  X"20",  X"60",  X"A0",  X"A0",  X"A0",
  X"20",  X"60",  X"40",  X"20",  X"40",  X"FF",  X"60",  X"20",
  X"40",  X"FF",  X"20",  X"FF",  X"20",  X"FF",  X"00",  X"60",
  X"80",  X"20",  X"60",  X"A0",  X"A0",  X"00",  X"60",  X"00",
  X"A0",  X"E0",  X"00",  X"80",  X"FF",  X"20",  X"E0",  X"FF",
  X"A0",  X"20",  X"00",  X"BF",  X"60",  X"80",  X"FF",  X"3F",
  X"60",  X"20",  X"00",  X"FF",  X"20",  X"FF",  X"60",  X"00",
  X"00",  X"20",  X"FF",  X"00",  X"A0",  X"60",  X"40",  X"FF",
  X"20",  X"FE",  X"A0",  X"A2",  X"40",  X"80",  X"00",  X"A2",
  X"E0",  X"FF",  X"00",  X"00",  X"80",  X"40",  X"A2",  X"A0",
  X"00",  X"00",  X"20",  X"40",  X"80",  X"70",  X"80",  X"00",
  X"6F",  X"40",  X"00",  X"00",  X"3F",  X"00",  X"20",  X"00",
  X"80",  X"A0",  X"A2",  X"40",  X"A2",  X"A0",  X"40",  X"00",
  X"60",  X"20",  X"00",  X"3F",  X"BF",  X"C0",  X"E0",  X"20",
  X"80",  X"E0",  X"20",  X"E0",  X"A0",  X"00",  X"E0",  X"00",
  X"A2",  X"40",  X"00",  X"A2",  X"00",  X"A2",  X"40",  X"FE",
  X"A2",  X"FE",  X"60",  X"FF",  X"60",  X"FE",  X"00",  X"65",
  X"20",  X"20",  X"FE",  X"20",  X"60",  X"FF",  X"20",  X"60",
  X"00",  X"61",  X"A0",  X"20",  X"FF",  X"20",  X"20",  X"20",
  X"80",  X"40",  X"60",  X"FF",  X"00",  X"23",  X"FE",  X"20",
  X"20",  X"20",  X"FE",  X"20",  X"20",  X"FE",  X"A0",  X"00",
  X"65",  X"A0",  X"20",  X"FE",  X"20",  X"AF",  X"FF",  X"E0",
  X"60",  X"40",  X"E0",  X"FF",  X"A0",  X"FF",  X"60",  X"E0",
  X"10",  X"00",  X"00",  X"FF",  X"62",  X"FF",  X"20",  X"23",
  X"FE",  X"20",  X"A0",  X"20",  X"FE",  X"20",  X"60",  X"40",
  X"FF",  X"60",  X"FF",  X"E0",  X"00",  X"20",  X"C0",  X"1F",
  X"40",  X"00",  X"00",  X"20",  X"C0",  X"1E",  X"40",  X"00",
  X"BF",  X"00",  X"00",  X"1C",  X"21",  X"3F",  X"00",  X"21",
  X"E0",  X"00",  X"60",  X"FF",  X"00",  X"00",  X"E0",  X"00",
  X"33",  X"24",  X"24",  X"31",  X"24",  X"24",  X"24",  X"24",
  X"24",  X"24",  X"30",  X"31",  X"24",  X"30",  X"32",  X"24",
  X"31",  X"31",  X"31",  X"31",  X"31",  X"31",  X"31",  X"31",
  X"31",  X"31",  X"24",  X"24",  X"24",  X"24",  X"24",  X"24",
  X"24",  X"24",  X"24",  X"30",  X"28",  X"33",  X"24",  X"33",
  X"24",  X"24",  X"24",  X"24",  X"33",  X"24",  X"24",  X"27",
  X"24",  X"24",  X"24",  X"32",  X"24",  X"27",  X"24",  X"24",
  X"33",  X"24",  X"24",  X"24",  X"24",  X"24",  X"24",  X"24",
  X"24",  X"24",  X"24",  X"30",  X"28",  X"33",  X"33",  X"33",
  X"32",  X"28",  X"24",  X"24",  X"31",  X"24",  X"30",  X"27",
  X"31",  X"31",  X"24",  X"32",  X"24",  X"27",  X"24",  X"24",
  X"31",  X"BF",  X"60",  X"60",  X"00",  X"00",  X"60",  X"E0",
  X"20",  X"10",  X"00",  X"60",  X"60",  X"E0",  X"00",  X"B8",
  X"11",  X"00",  X"00",  X"60",  X"A0",  X"62",  X"03",  X"B8",
  X"00",  X"62",  X"20",  X"00",  X"60",  X"20",  X"60",  X"03",
  X"00",  X"60",  X"60",  X"02",  X"00",  X"60",  X"A0",  X"02",
  X"60",  X"A0",  X"02",  X"60",  X"BF",  X"BF",  X"BF",  X"BF",
  X"B8",  X"B8",  X"B8",  X"B8",  X"00",  X"00",  X"A0",  X"60",
  X"20",  X"00",  X"80",  X"A0",  X"00",  X"80",  X"A0",  X"00",
  X"60",  X"00",  X"20",  X"00",  X"60",  X"00",  X"60",  X"FF",
  X"20",  X"00",  X"00",  X"00",  X"20",  X"00",  X"20",  X"BF",
  X"BF",  X"60",  X"80",  X"BF",  X"60",  X"02",  X"BF",  X"00",
  X"00",  X"00",  X"60",  X"60",  X"05",  X"A0",  X"BF",  X"3F",
  X"80",  X"60",  X"20",  X"20",  X"20",  X"20",  X"60",  X"A0",
  X"7F",  X"60",  X"00",  X"60",  X"60",  X"05",  X"20",  X"BD",
  X"BF",  X"B9",  X"B9",  X"20",  X"BD",  X"20",  X"20",  X"01",
  X"20",  X"B9",  X"A0",  X"B9",  X"01",  X"B9",  X"BF",  X"60",
  X"01",  X"20",  X"20",  X"20",  X"BF",  X"00",  X"BF",  X"BF",
  X"60",  X"A0",  X"BF",  X"BF",  X"60",  X"01",  X"20",  X"B9",
  X"60",  X"01",  X"B9",  X"B9",  X"80",  X"60",  X"00",  X"60",
  X"00",  X"B9",  X"00",  X"20",  X"00",  X"00",  X"00",  X"3F",
  X"20",  X"00",  X"00",  X"60",  X"40",  X"60",  X"BF",  X"BF",
  X"E0",  X"20",  X"BF",  X"E0",  X"FF",  X"BF",  X"B8",  X"00",
  X"FF",  X"BF",  X"20",  X"01",  X"B8",  X"3F",  X"20",  X"FF",
  X"00",  X"00",  X"00",  X"00",  X"20",  X"B9",  X"00",  X"BF",
  X"80",  X"BF",  X"BF",  X"60",  X"BF",  X"60",  X"00",  X"20",
  X"00",  X"FF",  X"BF",  X"20",  X"01",  X"00",  X"21",  X"01",
  X"60",  X"20",  X"00",  X"20",  X"BF",  X"40",  X"BF",  X"BF",
  X"60",  X"60",  X"02",  X"BF",  X"20",  X"00",  X"BF",  X"B9",
  X"00",  X"20",  X"00",  X"20",  X"00",  X"B9",  X"20",  X"00",
  X"BF",  X"3F",  X"20",  X"00",  X"20",  X"20",  X"00",  X"20",
  X"BF",  X"BF",  X"60",  X"A0",  X"BF",  X"60",  X"FF",  X"BF",
  X"00",  X"FF",  X"00",  X"20",  X"01",  X"3F",  X"20",  X"FF",
  X"00",  X"20",  X"B9",  X"00",  X"BF",  X"00",  X"BF",  X"60",
  X"BF",  X"60",  X"00",  X"BF",  X"00",  X"FE",  X"BF",  X"20",
  X"01",  X"A0",  X"BF",  X"B9",  X"00",  X"00",  X"00",  X"20",
  X"01",  X"00",  X"BF",  X"A0",  X"FF",  X"00",  X"A0",  X"0E",
  X"00",  X"FF",  X"80",  X"00",  X"A1",  X"80",  X"40",  X"00",
  X"FF",  X"00",  X"20",  X"20",  X"00",  X"C0",  X"20",  X"00",
  X"C0",  X"E0",  X"00",  X"E0",  X"20",  X"20",  X"BF",  X"A0",
  X"00",  X"3F",  X"BE",  X"A0",  X"00",  X"B8",  X"A0",  X"00",
  X"60",  X"60",  X"60",  X"03",  X"60",  X"03",  X"BE",  X"60",
  X"FF",  X"60",  X"60",  X"60",  X"FF",  X"C0",  X"B8",  X"20",
  X"00",  X"80",  X"60",  X"00",  X"20",  X"FF",  X"80",  X"00",
  X"C0",  X"00",  X"E0",  X"20",  X"FF",  X"20",  X"20",  X"20",
  X"00",  X"C0",  X"20",  X"00",  X"C0",  X"E0",  X"00",  X"E0",
  X"20",  X"FF",  X"20",  X"00",  X"E0",  X"20",  X"FF",  X"20",
  X"20",  X"20",  X"02",  X"20",  X"C0",  X"E0",  X"60",  X"03",
  X"00",  X"20",  X"FF",  X"20",  X"00",  X"BE",  X"20",  X"01",
  X"20",  X"BE",  X"20",  X"40",  X"00",  X"B9",  X"B9",  X"B9",
  X"20",  X"BF",  X"60",  X"FE",  X"20",  X"B9",  X"60",  X"B9",
  X"20",  X"FE",  X"B9",  X"B9",  X"00",  X"60",  X"FE",  X"60",
  X"00",  X"B9",  X"00",  X"20",  X"00",  X"00",  X"00",  X"3F",
  X"20",  X"00",  X"00",  X"60",  X"40",  X"60",  X"BF",  X"BF",
  X"E0",  X"20",  X"BF",  X"E0",  X"FF",  X"BF",  X"B8",  X"00",
  X"FE",  X"BF",  X"20",  X"00",  X"B8",  X"3F",  X"20",  X"FF",
  X"00",  X"00",  X"00",  X"00",  X"20",  X"B9",  X"00",  X"BF",
  X"80",  X"BF",  X"BF",  X"60",  X"BF",  X"60",  X"FE",  X"20",
  X"00",  X"FE",  X"BF",  X"20",  X"00",  X"BF",  X"60",  X"FE",
  X"00",  X"20",  X"FE",  X"B9",  X"BF",  X"20",  X"BF",  X"20",
  X"20",  X"BF",  X"00",  X"BF",  X"BF",  X"60",  X"A0",  X"BF",
  X"BF",  X"60",  X"FE",  X"20",  X"00",  X"FE",  X"BF",  X"20",
  X"00",  X"B9",  X"60",  X"FE",  X"00",  X"B9",  X"00",  X"60",
  X"FE",  X"60",  X"00",  X"B9",  X"00",  X"20",  X"00",  X"00",
  X"00",  X"3F",  X"20",  X"00",  X"00",  X"60",  X"40",  X"60",
  X"BF",  X"BF",  X"E0",  X"20",  X"BF",  X"E0",  X"FF",  X"BF",
  X"B8",  X"00",  X"FD",  X"BF",  X"20",  X"00",  X"B8",  X"3F",
  X"20",  X"FF",  X"00",  X"00",  X"00",  X"00",  X"20",  X"B9",
  X"00",  X"BF",  X"80",  X"BF",  X"BF",  X"60",  X"BF",  X"60",
  X"FE",  X"20",  X"00",  X"FD",  X"BF",  X"20",  X"00",  X"00",
  X"FE",  X"B9",  X"00",  X"B8",  X"00",  X"B8",  X"60",  X"40",
  X"8A",  X"00",  X"00",  X"BF",  X"20",  X"20",  X"00",  X"60",
  X"BF",  X"00",  X"BF",  X"60",  X"A0",  X"BF",  X"BF",  X"60",
  X"03",  X"20",  X"BF",  X"B8",  X"40",  X"00",  X"20",  X"20",
  X"FE",  X"20",  X"20",  X"20",  X"B8",  X"00",  X"BF",  X"BF",
  X"60",  X"A0",  X"BF",  X"BF",  X"60",  X"04",  X"20",  X"B8",
  X"7F",  X"60",  X"FE",  X"60",  X"02",  X"B9",  X"20",  X"00",
  X"BF",  X"7F",  X"60",  X"02",  X"20",  X"20",  X"00",  X"20",
  X"BF",  X"BF",  X"60",  X"A0",  X"BF",  X"60",  X"FF",  X"BF",
  X"00",  X"FD",  X"00",  X"20",  X"00",  X"00",  X"FF",  X"7F",
  X"00",  X"FD",  X"BF",  X"20",  X"FE",  X"BF",  X"A0",  X"00",
  X"60",  X"A0",  X"0D",  X"00",  X"60",  X"60",  X"60",  X"62",
  X"00",  X"00",  X"60",  X"00",  X"00",  X"E0",  X"00",  X"E0",
  X"3F",  X"06",  X"00",  X"20",  X"04",  X"60",  X"60",  X"00",
  X"E0",  X"A0",  X"FD",  X"BF",  X"60",  X"A0",  X"FD",  X"60",
  X"62",  X"00",  X"00",  X"FF",  X"60",  X"BE",  X"B9",  X"60",
  X"BE",  X"BE",  X"24",  X"BE",  X"BE",  X"BE",  X"BF",  X"BE",
  X"BE",  X"00",  X"1B",  X"BE",  X"00",  X"1C",  X"20",  X"00",
  X"BE",  X"1B",  X"00",  X"1B",  X"00",  X"A0",  X"BE",  X"00",
  X"00",  X"FD",  X"00",  X"20",  X"00",  X"BE",  X"0B",  X"00",
  X"20",  X"00",  X"3F",  X"BE",  X"60",  X"00",  X"00",  X"60",
  X"60",  X"60",  X"1B",  X"00",  X"E0",  X"00",  X"60",  X"01",
  X"20",  X"C0",  X"BF",  X"20",  X"BF",  X"20",  X"20",  X"BF",
  X"00",  X"BF",  X"BF",  X"60",  X"A0",  X"BF",  X"BF",  X"60",
  X"01",  X"20",  X"00",  X"B8",  X"A0",  X"80",  X"8A",  X"00",
  X"00",  X"B8",  X"B8",  X"BF",  X"20",  X"E0",  X"00",  X"BF",
  X"80",  X"BF",  X"BF",  X"60",  X"BF",  X"60",  X"01",  X"20",
  X"B8",  X"20",  X"BF",  X"B8",  X"00",  X"BF",  X"BF",  X"60",
  X"80",  X"BF",  X"BF",  X"60",  X"FD",  X"20",  X"00",  X"FC",
  X"BF",  X"20",  X"FF",  X"00",  X"FD",  X"20",  X"00",  X"FC",
  X"BF",  X"20",  X"FF",  X"00",  X"FD",  X"00",  X"1B",  X"60",
  X"FC",  X"00",  X"0C",  X"00",  X"FC",  X"60",  X"1B",  X"60",
  X"FF",  X"60",  X"60",  X"02",  X"B8",  X"40",  X"01",  X"20",
  X"20",  X"B8",  X"00",  X"BF",  X"BF",  X"60",  X"80",  X"BF",
  X"BF",  X"60",  X"02",  X"20",  X"BF",  X"B8",  X"40",  X"60",
  X"02",  X"60",  X"01",  X"B9",  X"20",  X"00",  X"BF",  X"7F",
  X"60",  X"01",  X"20",  X"20",  X"00",  X"20",  X"BF",  X"BF",
  X"60",  X"A0",  X"BF",  X"60",  X"FF",  X"BF",  X"00",  X"FC",
  X"00",  X"20",  X"FF",  X"00",  X"FF",  X"7F",  X"BE",  X"BE",
  X"FE",  X"20",  X"FF",  X"60",  X"FF",  X"60",  X"01",  X"B9",
  X"20",  X"00",  X"BF",  X"7F",  X"60",  X"01",  X"20",  X"20",
  X"00",  X"20",  X"BF",  X"BF",  X"60",  X"A0",  X"BF",  X"60",
  X"FF",  X"BF",  X"00",  X"FC",  X"00",  X"20",  X"FF",  X"00",
  X"FF",  X"7F",  X"FD",  X"C0",  X"E0",  X"FD",  X"E0",  X"1B",
  X"60",  X"60",  X"FF",  X"60",  X"C0",  X"20",  X"00",  X"E0",
  X"00",  X"80",  X"20",  X"FC",  X"60",  X"60",  X"01",  X"20",
  X"01",  X"BF",  X"C0",  X"20",  X"E0",  X"BD",  X"BD",  X"00",
  X"BF",  X"60",  X"B9",  X"40",  X"20",  X"FC",  X"B9",  X"20",
  X"00",  X"C0",  X"20",  X"00",  X"00",  X"E0",  X"FC",  X"40",
  X"80",  X"20",  X"FC",  X"60",  X"80",  X"FC",  X"60",  X"BF",
  X"80",  X"FC",  X"60",  X"80",  X"20",  X"FC",  X"60",  X"7F",
  X"20",  X"80",  X"20",  X"20",  X"00",  X"40",  X"7F",  X"60",
  X"FF",  X"A0",  X"FC",  X"7F",  X"C0",  X"00",  X"00",  X"E0",
  X"E0",  X"20",  X"20",  X"B8",  X"20",  X"FD",  X"20",  X"80",
  X"20",  X"FC",  X"60",  X"80",  X"60",  X"60",  X"60",  X"02",
  X"A0",  X"FC",  X"20",  X"00",  X"60",  X"20",  X"00",  X"B8",
  X"20",  X"00",  X"C0",  X"E0",  X"E0",  X"00",  X"20",  X"A0",
  X"FD",  X"20",  X"20",  X"FD",  X"BF",  X"20",  X"FD",  X"20",
  X"80",  X"60",  X"03",  X"A0",  X"7F",  X"20",  X"60",  X"FC",
  X"20",  X"80",  X"A0",  X"A0",  X"80",  X"80",  X"7F",  X"60",
  X"FF",  X"A0",  X"A0",  X"FC",  X"3F",  X"FC",  X"7F",  X"80",
  X"20",  X"FC",  X"60",  X"BF",  X"C0",  X"E0",  X"02",  X"E0",
  X"60",  X"00",  X"20",  X"00",  X"BF",  X"A0",  X"01",  X"00",
  X"20",  X"0E",  X"00",  X"20",  X"00",  X"B9",  X"00",  X"40",
  X"02",  X"00",  X"B9",  X"00",  X"B9",  X"FD",  X"20",  X"00",
  X"E0",  X"20",  X"FF",  X"B8",  X"C0",  X"FF",  X"E0",  X"BF",
  X"60",  X"FF",  X"80",  X"BF",  X"80",  X"FC",  X"60",  X"80",
  X"20",  X"FC",  X"60",  X"BF",  X"01",  X"60",  X"01",  X"60",
  X"01",  X"A0",  X"20",  X"00",  X"00",  X"BF",  X"0E",  X"20",
  X"BF",  X"B8",  X"B9",  X"E0",  X"14",  X"B8",  X"20",  X"01",
  X"00",  X"B8",  X"60",  X"40",  X"8A",  X"00",  X"00",  X"20",
  X"20",  X"00",  X"B9",  X"20",  X"B9",  X"E0",  X"FD",  X"20",
  X"E0",  X"FB",  X"40",  X"B8",  X"60",  X"80",  X"FF",  X"60",
  X"60",  X"FF",  X"C0",  X"B8",  X"FD",  X"40",  X"60",  X"00",
  X"BE",  X"00",  X"00",  X"20",  X"16",  X"FF",  X"20",  X"20",
  X"00",  X"16",  X"C0",  X"20",  X"FF",  X"00",  X"00",  X"60",
  X"B8",  X"BF",  X"BF",  X"FC",  X"C0",  X"FE",  X"C0",  X"20",
  X"20",  X"00",  X"20",  X"BF",  X"BF",  X"60",  X"A0",  X"BF",
  X"60",  X"FE",  X"BF",  X"00",  X"FB",  X"BF",  X"20",  X"FD",
  X"00",  X"FE",  X"B8",  X"00",  X"FB",  X"BF",  X"20",  X"FD",
  X"00",  X"FE",  X"00",  X"20",  X"B9",  X"00",  X"BF",  X"40",
  X"BF",  X"60",  X"BF",  X"BF",  X"60",  X"FE",  X"20",  X"FF",
  X"00",  X"BF",  X"20",  X"20",  X"0E",  X"00",  X"C0",  X"A0",
  X"00",  X"BD",  X"02",  X"00",  X"3F",  X"02",  X"00",  X"FE",
  X"E0",  X"20",  X"00",  X"BF",  X"00",  X"20",  X"FC",  X"20",
  X"20",  X"B9",  X"00",  X"BF",  X"40",  X"20",  X"FC",  X"BF",
  X"BF",  X"0D",  X"20",  X"BF",  X"B8",  X"E0",  X"FF",  X"B9",
  X"BF",  X"20",  X"BF",  X"0E",  X"20",  X"A0",  X"01",  X"20",
  X"20",  X"B9",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"BF",  X"40",  X"A0",  X"01",  X"A0",  X"BD",  X"02",
  X"BF",  X"3F",  X"01",  X"60",  X"00",  X"40",  X"01",  X"40",
  X"FF",  X"A0",  X"00",  X"00",  X"B9",  X"60",  X"01",  X"20",
  X"B9",  X"FC",  X"B9",  X"00",  X"20",  X"BF",  X"80",  X"BF",
  X"BF",  X"60",  X"60",  X"00",  X"BF",  X"20",  X"BF",  X"20",
  X"00",  X"60",  X"BF",  X"00",  X"BF",  X"60",  X"A0",  X"BF",
  X"BF",  X"60",  X"00",  X"20",  X"BF",  X"B8",  X"C0",  X"20",
  X"C0",  X"00",  X"BF",  X"80",  X"BF",  X"FD",  X"60",  X"20",
  X"B9",  X"00",  X"BF",  X"40",  X"BF",  X"60",  X"BF",  X"BF",
  X"60",  X"00",  X"20",  X"00",  X"FA",  X"BF",  X"20",  X"FD",
  X"00",  X"20",  X"FB",  X"20",  X"20",  X"20",  X"00",  X"60",
  X"BF",  X"00",  X"BF",  X"60",  X"FD",  X"A0",  X"A0",  X"FE",
  X"20",  X"FE",  X"20",  X"00",  X"FA",  X"BF",  X"20",  X"FD",
  X"00",  X"FC",  X"BF",  X"20",  X"00",  X"BF",  X"B9",  X"20",
  X"E0",  X"B9",  X"FC",  X"20",  X"20",  X"20",  X"00",  X"60",
  X"BF",  X"00",  X"BF",  X"60",  X"A0",  X"BF",  X"BF",  X"60",
  X"00",  X"20",  X"BF",  X"60",  X"00",  X"B8",  X"20",  X"20",
  X"B8",  X"00",  X"BF",  X"BF",  X"A0",  X"E0",  X"BF",  X"BF",
  X"A0",  X"01",  X"20",  X"BF",  X"00",  X"60",  X"00",  X"60",
  X"00",  X"B9",  X"20",  X"00",  X"BF",  X"7F",  X"60",  X"00",
  X"60",  X"60",  X"40",  X"60",  X"BF",  X"BF",  X"A0",  X"E0",
  X"BF",  X"A0",  X"FF",  X"BF",  X"00",  X"FA",  X"00",  X"20",
  X"FC",  X"00",  X"FF",  X"7F",  X"E0",  X"FB",  X"20",  X"FF",
  X"20",  X"00",  X"FA",  X"BF",  X"20",  X"FC",  X"00",  X"FD",
  X"BF",  X"00",  X"FA",  X"BF",  X"20",  X"FC",  X"00",  X"FF",
  X"BF",  X"00",  X"FA",  X"BF",  X"20",  X"FC",  X"00",  X"FF",
  X"20",  X"00",  X"FA",  X"BF",  X"20",  X"FC",  X"00",  X"FF",
  X"BF",  X"B9",  X"13",  X"20",  X"00",  X"00",  X"60",  X"00",
  X"FB",  X"B9",  X"BF",  X"60",  X"00",  X"00",  X"BF",  X"FC",
  X"60",  X"FA",  X"BF",  X"20",  X"FC",  X"60",  X"BF",  X"FC",
  X"60",  X"FE",  X"20",  X"80",  X"20",  X"FA",  X"60",  X"12",
  X"B8",  X"20",  X"00",  X"20",  X"21",  X"60",  X"00",  X"00",
  X"20",  X"60",  X"01",  X"60",  X"00",  X"20",  X"B8",  X"BF",
  X"B9",  X"BF",  X"60",  X"01",  X"00",  X"BF",  X"A0",  X"A0",
  X"B9",  X"BF",  X"B9",  X"A0",  X"00",  X"03",  X"BF",  X"60",
  X"00",  X"00",  X"60",  X"00",  X"20",  X"00",  X"60",  X"C0",
  X"01",  X"60",  X"40",  X"B9",  X"8A",  X"00",  X"00",  X"BF",
  X"BF",  X"60",  X"80",  X"00",  X"3F",  X"60",  X"00",  X"B8",
  X"60",  X"00",  X"60",  X"BF",  X"7F",  X"00",  X"60",  X"80",
  X"00",  X"B8",  X"60",  X"20",  X"00",  X"20",  X"20",  X"20",
  X"7F",  X"BF",  X"60",  X"01",  X"BF",  X"20",  X"BF",  X"60",
  X"00",  X"BF",  X"60",  X"20",  X"BF",  X"BF",  X"BF",  X"B8",
  X"60",  X"BF",  X"80",  X"B8",  X"B8",  X"00",  X"40",  X"60",
  X"B9",  X"A0",  X"00",  X"00",  X"20",  X"B9",  X"BF",  X"20",
  X"00",  X"60",  X"40",  X"60",  X"FB",  X"B9",  X"20",  X"FF",
  X"B9",  X"FF",  X"60",  X"00",  X"F9",  X"BF",  X"20",  X"FC",
  X"00",  X"FB",  X"B8",  X"B9",  X"60",  X"20",  X"40",  X"FB",
  X"B9",  X"60",  X"B9",  X"40",  X"BF",  X"80",  X"BF",  X"A0",
  X"BF",  X"BF",  X"A0",  X"00",  X"60",  X"00",  X"F9",  X"BF",
  X"20",  X"FC",  X"00",  X"B8",  X"60",  X"40",  X"60",  X"BF",
  X"BF",  X"60",  X"80",  X"BF",  X"60",  X"FA",  X"BF",  X"FC",
  X"00",  X"20",  X"00",  X"B9",  X"20",  X"E0",  X"B9",  X"F9",
  X"20",  X"00",  X"B9",  X"20",  X"B9",  X"E0",  X"FA",  X"20",
  X"A0",  X"F7",  X"60",  X"20",  X"00",  X"20",  X"20",  X"0C",
  X"BF",  X"A0",  X"00",  X"BF",  X"BF",  X"00",  X"00",  X"40",
  X"00",  X"00",  X"80",  X"00",  X"60",  X"B9",  X"40",  X"FA",
  X"B9",  X"62",  X"FB",  X"60",  X"17",  X"3F",  X"E0",  X"00",
  X"00",  X"00",  X"00",  X"FE",  X"B9",  X"00",  X"60",  X"00",
  X"BF",  X"B8",  X"C0",  X"00",  X"60",  X"20",  X"FF",  X"20",
  X"FF",  X"60",  X"20",  X"FF",  X"00",  X"FF",  X"BF",  X"80",
  X"00",  X"00",  X"20",  X"40",  X"60",  X"80",  X"FF",  X"BF",
  X"FF",  X"60",  X"A0",  X"20",  X"BF",  X"20",  X"00",  X"BF",
  X"3F",  X"00",  X"00",  X"FE",  X"BF",  X"00",  X"F9",  X"BF",
  X"20",  X"FB",  X"00",  X"FE",  X"BF",  X"60",  X"A0",  X"00",
  X"FB",  X"60",  X"A0",  X"FF",  X"20",  X"00",  X"B8",  X"00",
  X"20",  X"14",  X"BF",  X"20",  X"20",  X"00",  X"13",  X"80",
  X"B8",  X"20",  X"FF",  X"00",  X"20",  X"BF",  X"00",  X"BF",
  X"40",  X"00",  X"BF",  X"FF",  X"B8",  X"C0",  X"E0",  X"80",
  X"40",  X"FF",  X"A0",  X"FF",  X"B8",  X"BF",  X"FF",  X"00",
  X"00",  X"00",  X"20",  X"B9",  X"FE",  X"B9",  X"C0",  X"60",
  X"00",  X"00",  X"BF",  X"80",  X"FE",  X"60",  X"20",  X"00",
  X"40",  X"20",  X"B8",  X"40",  X"FF",  X"20",  X"00",  X"B9",
  X"E0",  X"C0",  X"8A",  X"00",  X"00",  X"00",  X"20",  X"C0",
  X"BF",  X"FE",  X"80",  X"20",  X"00",  X"FE",  X"BF",  X"BF",
  X"FE",  X"80",  X"C0",  X"A0",  X"FC",  X"E0",  X"80",  X"60",
  X"F9",  X"3F",  X"60",  X"00",  X"A0",  X"00",  X"60",  X"20",
  X"FE",  X"B9",  X"60",  X"20",  X"FE",  X"40",  X"00",  X"A0",
  X"20",  X"FE",  X"20",  X"A0",  X"FE",  X"20",  X"FE",  X"00",
  X"60",  X"60",  X"FB",  X"60",  X"00",  X"00",  X"62",  X"00",
  X"00",  X"00",  X"00",  X"C0",  X"F8",  X"40",  X"00",  X"BF",
  X"60",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"3F",  X"00",  X"00",  X"C0",  X"20",  X"00",  X"E0",  X"00",
  X"00",  X"BF",  X"20",  X"00",  X"00",  X"FF",  X"3F",  X"00",
  X"00",  X"62",  X"00",  X"00",  X"00",  X"00",  X"C0",  X"FF",
  X"40",  X"00",  X"BF",  X"60",  X"00",  X"00",  X"E0",  X"00",
  X"80",  X"C0",  X"BF",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"FF",  X"00",  X"3F",  X"00",  X"20",  X"C0",  X"40",  X"00",
  X"20",  X"00",  X"00",  X"20",  X"60",  X"00",  X"00",  X"20",
  X"00",  X"20",  X"40",  X"80",  X"60",  X"00",  X"FF",  X"40",
  X"80",  X"80",  X"60",  X"80",  X"C0",  X"60",  X"00",  X"00",
  X"00",  X"E0",  X"C0",  X"00",  X"20",  X"00",  X"00",  X"FF",
  X"00",  X"3F",  X"FF",  X"C0",  X"20",  X"00",  X"00",  X"E0",
  X"3F",  X"00",  X"E0",  X"00",  X"20",  X"E0",  X"00",  X"60",
  X"00",  X"80",  X"00",  X"E0",  X"3F",  X"80",  X"FF",  X"3F",
  X"00",  X"00",  X"00",  X"62",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"C0",  X"FF",  X"40",  X"00",  X"BF",  X"00",  X"11",
  X"21",  X"20",  X"00",  X"21",  X"00",  X"11",  X"60",  X"20",
  X"00",  X"60",  X"00",  X"A0",  X"00",  X"40",  X"BF",  X"67",
  X"00",  X"A0",  X"A7",  X"7F",  X"A0",  X"BF",  X"60",  X"40",
  X"E0",  X"20",  X"21",  X"00",  X"11",  X"60",  X"20",  X"00",
  X"60",  X"00",  X"A0",  X"60",  X"00",  X"60",  X"40",  X"E0",
  X"20",  X"60",  X"FF",  X"40",  X"E0",  X"20",  X"B8",  X"00",
  X"63",  X"80",  X"00",  X"FF",  X"07",  X"80",  X"63",  X"80",
  X"00",  X"A0",  X"A0",  X"3F",  X"E0",  X"A0",  X"FF",  X"A0",
  X"AF",  X"BF",  X"60",  X"7F",  X"60",  X"40",  X"60",  X"60",
  X"E0",  X"20",  X"F8",  X"F7",  X"80",  X"63",  X"80",  X"00",
  X"A0",  X"A0",  X"7F",  X"20",  X"A0",  X"3F",  X"E0",  X"A0",
  X"FF",  X"A0",  X"AF",  X"BF",  X"60",  X"7F",  X"60",  X"40",
  X"60",  X"60",  X"60",  X"E0",  X"20",  X"E0",  X"E0",  X"00",
  X"60",  X"BF",  X"60",  X"60",  X"00",  X"00",  X"BF",  X"E0",
  X"E0",  X"00",  X"3F",  X"60",  X"40",  X"E0",  X"20",  X"21",
  X"00",  X"10",  X"60",  X"20",  X"00",  X"60",  X"FF",  X"A0",
  X"60",  X"FF",  X"40",  X"60",  X"A0",  X"A0",  X"00",  X"A0",
  X"E0",  X"3F",  X"21",  X"00",  X"10",  X"60",  X"20",  X"FF",
  X"60",  X"00",  X"20",  X"A0",  X"60",  X"00",  X"00",  X"C0",
  X"60",  X"00",  X"20",  X"C0",  X"40",  X"20",  X"20",  X"60",
  X"20",  X"60",  X"60",  X"40",  X"E0",  X"00",  X"FF",  X"80",
  X"67",  X"FF",  X"A0",  X"A0",  X"FF",  X"A0",  X"AF",  X"BF",
  X"60",  X"7F",  X"60",  X"40",  X"60",  X"E0",  X"20",  X"60",
  X"60",  X"FF",  X"BF",  X"E0",  X"3F",  X"A0",  X"A0",  X"3F",
  X"60",  X"A0",  X"7F",  X"20",  X"A0",  X"3F",  X"E0",  X"A0",
  X"FF",  X"A0",  X"AF",  X"BF",  X"60",  X"7F",  X"60",  X"40",
  X"60",  X"60",  X"60",  X"60",  X"E0",  X"20",  X"7F",  X"60",
  X"60",  X"FF",  X"3F",  X"BF",  X"60",  X"60",  X"00",  X"00",
  X"C0",  X"60",  X"00",  X"20",  X"20",  X"C0",  X"20",  X"40",
  X"20",  X"20",  X"60",  X"20",  X"60",  X"60",  X"60",  X"40",
  X"E0",  X"00",  X"A0",  X"A0",  X"FF",  X"3F",  X"60",  X"40",
  X"E0",  X"20",  X"BF",  X"00",  X"62",  X"20",  X"00",  X"00",
  X"20",  X"60",  X"00",  X"00",  X"20",  X"60",  X"A0",  X"A0",
  X"00",  X"00",  X"20",  X"A0",  X"00",  X"00",  X"20",  X"60",
  X"00",  X"60",  X"00",  X"20",  X"20",  X"20",  X"E0",  X"00",
  X"20",  X"20",  X"E0",  X"20",  X"20",  X"00",  X"20",  X"20",
  X"E0",  X"20",  X"06",  X"00",  X"FF",  X"20",  X"09",  X"00",
  X"FF",  X"20",  X"A0",  X"FF",  X"3F",  X"A0",  X"00",  X"20",
  X"E0",  X"20",  X"FF",  X"20",  X"60",  X"00",  X"7F",  X"20",
  X"40",  X"00",  X"20",  X"06",  X"62",  X"20",  X"20",  X"7F",
  X"20",  X"20",  X"20",  X"E0",  X"00",  X"FF",  X"20",  X"BF",
  X"20",  X"60",  X"00",  X"C0",  X"00",  X"20",  X"E0",  X"60",
  X"00",  X"40",  X"60",  X"60",  X"60",  X"00",  X"11",  X"FF",
  X"60",  X"20",  X"60",  X"00",  X"20",  X"00",  X"00",  X"63",
  X"00",  X"20",  X"20",  X"00",  X"C0",  X"11",  X"00",  X"E0",
  X"80",  X"11",  X"00",  X"80",  X"60",  X"40",  X"C0",  X"80",
  X"A0",  X"C0",  X"80",  X"A0",  X"80",  X"C0",  X"C0",  X"A0",
  X"20",  X"80",  X"40",  X"A0",  X"A0",  X"FF",  X"E0",  X"A0",
  X"00",  X"00",  X"E0",  X"A0",  X"00",  X"00",  X"00",  X"20",
  X"00",  X"A0",  X"00",  X"7F",  X"00",  X"20",  X"40",  X"A0",
  X"00",  X"7F",  X"00",  X"FF",  X"FF",  X"20",  X"00",  X"0A",
  X"00",  X"20",  X"00",  X"00",  X"20",  X"E3",  X"00",  X"20",
  X"40",  X"40",  X"60",  X"20",  X"00",  X"C0",  X"40",  X"C0",
  X"C0",  X"E0",  X"80",  X"60",  X"60",  X"40",  X"40",  X"60",
  X"FF",  X"A0",  X"E0",  X"A0",  X"00",  X"60",  X"E0",  X"00",
  X"00",  X"00",  X"20",  X"00",  X"A0",  X"00",  X"7F",  X"20",
  X"E0",  X"00",  X"40",  X"A0",  X"00",  X"20",  X"7F",  X"00",
  X"FF",  X"FF",  X"20",  X"E0",  X"00",  X"BF",  X"20",  X"BF",
  X"BF",  X"60",  X"A0",  X"A0",  X"00",  X"BF",  X"20",  X"60",
  X"20",  X"BF",  X"20",  X"C0",  X"60",  X"BF",  X"00",  X"09",
  X"00",  X"BF",  X"20",  X"BF",  X"BF",  X"BF",  X"A0",  X"00",
  X"20",  X"40",  X"FC",  X"80",  X"80",  X"00",  X"00",  X"00",
  X"60",  X"00",  X"8A",  X"00",  X"00",  X"20",  X"40",  X"00",
  X"20",  X"00",  X"20",  X"00",  X"20",  X"00",  X"E0",  X"3F",
  X"A0",  X"40",  X"BF",  X"00",  X"09",  X"00",  X"80",  X"20",
  X"00",  X"BF",  X"A0",  X"00",  X"40",  X"00",  X"E0",  X"00",
  X"BF",  X"00",  X"63",  X"40",  X"BF",  X"A0",  X"00",  X"FC",
  X"00",  X"20",  X"20",  X"00",  X"00",  X"20",  X"60",  X"00",
  X"20",  X"20",  X"00",  X"E0",  X"00",  X"40",  X"00",  X"80",
  X"BF",  X"FF",  X"BF",  X"BF",  X"BF",  X"BF",  X"BF",  X"BF",
  X"00",  X"BF",  X"BF",  X"00",  X"00",  X"0A",  X"BF",  X"A0",
  X"00",  X"27",  X"BF",  X"BF",  X"BF",  X"00",  X"BF",  X"BF",
  X"BF",  X"BF",  X"40",  X"E4",  X"00",  X"20",  X"BF",  X"00",
  X"40",  X"E4",  X"00",  X"40",  X"80",  X"80",  X"BF",  X"A0",
  X"BF",  X"03",  X"19",  X"BF",  X"3B",  X"BF",  X"00",  X"84",
  X"00",  X"40",  X"20",  X"BF",  X"BF",  X"BF",  X"00",  X"60",
  X"00",  X"BF",  X"08",  X"A0",  X"89",  X"BF",  X"19",  X"00",
  X"A1",  X"88",  X"00",  X"A1",  X"09",  X"88",  X"60",  X"0A",
  X"1A",  X"BF",  X"00",  X"00",  X"BF",  X"19",  X"8A",  X"00",
  X"00",  X"FF",  X"20",  X"E0",  X"00",  X"BF",  X"E0",  X"00",
  X"E1",  X"C0",  X"8A",  X"00",  X"00",  X"BF",  X"FF",  X"7F",
  X"20",  X"40",  X"60",  X"00",  X"00",  X"00",  X"20",  X"E0",
  X"01",  X"00",  X"BF",  X"BF",  X"80",  X"E0",  X"00",  X"3F",
  X"E0",  X"00",  X"20",  X"FF",  X"20",  X"E0",  X"00",  X"20",
  X"01",  X"E0",  X"E0",  X"03",  X"E0",  X"01",  X"3F",  X"20",
  X"C0",  X"60",  X"20",  X"03",  X"BF",  X"20",  X"20",  X"20",
  X"03",  X"20",  X"00",  X"60",  X"60",  X"C0",  X"FF",  X"A0",
  X"A0",  X"20",  X"20",  X"BF",  X"40",  X"BF",  X"BF",  X"BF",
  X"0A",  X"00",  X"20",  X"00",  X"A0",  X"BF",  X"BF",  X"BF",
  X"00",  X"BF",  X"E0",  X"00",  X"BF",  X"60",  X"00",  X"00",
  X"E0",  X"A0",  X"A1",  X"02",  X"80",  X"09",  X"A0",  X"60",
  X"1A",  X"BF",  X"19",  X"89",  X"08",  X"BF",  X"20",  X"00",
  X"40",  X"00",  X"61",  X"09",  X"60",  X"0A",  X"00",  X"00",
  X"20",  X"61",  X"00",  X"60",  X"C0",  X"09",  X"40",  X"0A",
  X"00",  X"FF",  X"BF",  X"09",  X"60",  X"80",  X"1A",  X"BF",
  X"19",  X"89",  X"08",  X"BF",  X"20",  X"80",  X"FF",  X"A0",
  X"08",  X"0A",  X"00",  X"02",  X"BF",  X"0A",  X"00",  X"FE",
  X"BF",  X"BF",  X"BF",  X"60",  X"02",  X"BF",  X"FE",  X"BF",
  X"00",  X"80",  X"FF",  X"20",  X"FF",  X"00",  X"BF",  X"FC",
  X"3C",  X"BF",  X"BF",  X"00",  X"00",  X"FC",  X"80",  X"40",
  X"FF",  X"BF",  X"BF",  X"20",  X"20",  X"20",  X"3F",  X"20",
  X"20",  X"20",  X"BF",  X"BF",  X"BF",  X"BF",  X"09",  X"00",
  X"20",  X"00",  X"A0",  X"BF",  X"BF",  X"BF",  X"FF",  X"BF",
  X"E0",  X"02",  X"E0",  X"60",  X"00",  X"00",  X"A1",  X"00",
  X"80",  X"E0",  X"60",  X"01",  X"20",  X"60",  X"00",  X"09",
  X"00",  X"A2",  X"60",  X"00",  X"60",  X"80",  X"09",  X"E0",
  X"60",  X"FF",  X"A0",  X"09",  X"BF",  X"60",  X"00",  X"BF",
  X"00",  X"61",  X"0A",  X"00",  X"00",  X"00",  X"A0",  X"00",
  X"BF",  X"A0",  X"01",  X"E0",  X"BF",  X"00",  X"61",  X"09",
  X"00",  X"BF",  X"19",  X"09",  X"61",  X"88",  X"BF",  X"30",
  X"BF",  X"40",  X"FF",  X"01",  X"BF",  X"BF",  X"00",  X"A0",
  X"BF",  X"19",  X"89",  X"61",  X"88",  X"BF",  X"30",  X"BF",
  X"01",  X"40",  X"BF",  X"00",  X"61",  X"08",  X"BF",  X"0A",
  X"00",  X"01",  X"BF",  X"00",  X"0A",  X"00",  X"01",  X"00",
  X"BF",  X"20",  X"00",  X"BF",  X"00",  X"01",  X"20",  X"E0",
  X"01",  X"E0",  X"BF",  X"BF",  X"BF",  X"A0",  X"00",  X"BF",
  X"20",  X"00",  X"80",  X"00",  X"00",  X"00",  X"BF",  X"40",
  X"BF",  X"80",  X"40",  X"BF",  X"60",  X"00",  X"E0",  X"02",
  X"60",  X"00",  X"BF",  X"BF",  X"BF",  X"00",  X"0B",  X"00",
  X"BF",  X"00",  X"00",  X"0A",  X"BF",  X"00",  X"00",  X"07",
  X"00",  X"BF",  X"BF",  X"00",  X"BF",  X"80",  X"02",  X"00",
  X"BF",  X"BF",  X"00",  X"0A",  X"20",  X"BF",  X"00",  X"E0",
  X"BF",  X"00",  X"BF",  X"00",  X"00",  X"0A",  X"00",  X"BF",
  X"BF",  X"00",  X"E0",  X"01",  X"BF",  X"BF",  X"BF",  X"60",
  X"01",  X"20",  X"40",  X"60",  X"01",  X"20",  X"BF",  X"C0",
  X"BF",  X"80",  X"40",  X"60",  X"00",  X"00",  X"BF",  X"BF",
  X"00",  X"09",  X"00",  X"BF",  X"BF",  X"00",  X"A0",  X"00",
  X"00",  X"BF",  X"BF",  X"00",  X"09",  X"00",  X"BF",  X"BF",
  X"00",  X"BF",  X"20",  X"01",  X"BF",  X"A0",  X"02",  X"E0",
  X"E0",  X"00",  X"00",  X"20",  X"BF",  X"20",  X"00",  X"BF",
  X"BF",  X"BF",  X"00",  X"09",  X"00",  X"BF",  X"BF",  X"BF",
  X"BF",  X"60",  X"02",  X"BF",  X"BF",  X"BF",  X"00",  X"20",
  X"BF",  X"E0",  X"00",  X"FD",  X"00",  X"20",  X"00",  X"BF",
  X"07",  X"00",  X"00",  X"BF",  X"00",  X"09",  X"00",  X"20",
  X"A0",  X"00",  X"01",  X"20",  X"BF",  X"00",  X"07",  X"00",
  X"BF",  X"A0",  X"00",  X"BF",  X"E0",  X"00",  X"60",  X"60",
  X"02",  X"BF",  X"60",  X"01",  X"60",  X"00",  X"A0",  X"E0",
  X"00",  X"A0",  X"60",  X"01",  X"A0",  X"02",  X"BF",  X"80",
  X"80",  X"00",  X"A0",  X"00",  X"00",  X"20",  X"0A",  X"20",
  X"00",  X"01",  X"00",  X"00",  X"20",  X"20",  X"0A",  X"00",
  X"00",  X"00",  X"20",  X"00",  X"20",  X"0A",  X"A0",  X"FF",
  X"00",  X"40",  X"BF",  X"FE",  X"BF",  X"00",  X"A2",  X"89",
  X"60",  X"FE",  X"20",  X"01",  X"3F",  X"20",  X"20",  X"BF",
  X"3F",  X"FE",  X"20",  X"00",  X"20",  X"20",  X"0A",  X"E0",
  X"00",  X"00",  X"FC",  X"00",  X"20",  X"BF",  X"C0",  X"80",
  X"00",  X"FF",  X"A0",  X"BF",  X"20",  X"00",  X"20",  X"09",
  X"00",  X"00",  X"07",  X"00",  X"20",  X"00",  X"BF",  X"01",
  X"BF",  X"60",  X"BF",  X"01",  X"BF",  X"40",  X"FF",  X"00",
  X"20",  X"40",  X"E0",  X"00",  X"06",  X"00",  X"E0",  X"FE",
  X"00",  X"00",  X"20",  X"00",  X"00",  X"06",  X"00",  X"00",
  X"BF",  X"06",  X"00",  X"FD",  X"00",  X"01",  X"BF",  X"BF",
  X"40",  X"00",  X"40",  X"BF",  X"40",  X"40",  X"C0",  X"BF",
  X"BF",  X"20",  X"40",  X"BF",  X"A0",  X"00",  X"20",  X"BF",
  X"00",  X"BF",  X"BF",  X"80",  X"40",  X"00",  X"09",  X"20",
  X"BF",  X"BF",  X"FE",  X"BF",  X"BF",  X"00",  X"E0",  X"00",
  X"1A",  X"BF",  X"60",  X"00",  X"E1",  X"C0",  X"00",  X"61",
  X"89",  X"1A",  X"BF",  X"19",  X"08",  X"BF",  X"E0",  X"40",
  X"BF",  X"BF",  X"88",  X"0A",  X"00",  X"FD",  X"60",  X"00",
  X"21",  X"88",  X"0A",  X"00",  X"00",  X"A0",  X"00",  X"00",
  X"21",  X"61",  X"00",  X"20",  X"00",  X"88",  X"8A",  X"00",
  X"00",  X"BF",  X"00",  X"00",  X"09",  X"1A",  X"BF",  X"19",
  X"08",  X"09",  X"60",  X"0A",  X"40",  X"BF",  X"20",  X"80",
  X"00",  X"FF",  X"A0",  X"FC",  X"00",  X"BF",  X"20",  X"FE",
  X"BF",  X"BF",  X"FC",  X"BF",  X"40",  X"FE",  X"BF",  X"FC",
  X"40",  X"FE",  X"BF",  X"20",  X"60",  X"A0",  X"FE",  X"BF",
  X"BF",  X"60",  X"BF",  X"FC",  X"BF",  X"40",  X"FF",  X"00",
  X"20",  X"E0",  X"40",  X"20",  X"FC",  X"00",  X"00",  X"FD",
  X"00",  X"00",  X"BF",  X"06",  X"00",  X"BF",  X"FE",  X"00",
  X"20",  X"FD",  X"09",  X"A0",  X"FE",  X"00",  X"61",  X"09",
  X"0A",  X"00",  X"FE",  X"BF",  X"20",  X"BF",  X"20",  X"E0",
  X"40",  X"60",  X"FF",  X"20",  X"20",  X"80",  X"60",  X"01",
  X"BF",  X"7F",  X"80",  X"80",  X"40",  X"FE",  X"BF",  X"00",
  X"00",  X"20",  X"20",  X"09",  X"A0",  X"00",  X"FE",  X"00",
  X"00",  X"00",  X"00",  X"FD",  X"20",  X"60",  X"00",  X"A0",
  X"E1",  X"C0",  X"60",  X"89",  X"60",  X"FD",  X"20",  X"00",
  X"A2",  X"60",  X"00",  X"60",  X"80",  X"09",  X"E0",  X"60",
  X"FF",  X"A0",  X"FD",  X"BF",  X"BF",  X"19",  X"08",  X"A0",
  X"60",  X"BF",  X"E0",  X"00",  X"E1",  X"40",  X"BF",  X"BF",
  X"60",  X"C0",  X"BF",  X"00",  X"09",  X"00",  X"61",  X"20",
  X"09",  X"1A",  X"BF",  X"19",  X"BF",  X"20",  X"40",  X"60",
  X"40",  X"FF",  X"08",  X"7F",  X"80",  X"00",  X"61",  X"08",
  X"0A",  X"00",  X"FF",  X"BF",  X"08",  X"0A",  X"00",  X"FF",
  X"00",  X"00",  X"BF",  X"00",  X"BF",  X"60",  X"FF",  X"BF",
  X"FC",  X"00",  X"00",  X"A0",  X"FC",  X"08",  X"20",  X"20",
  X"00",  X"00",  X"BF",  X"FC",  X"00",  X"FF",  X"20",  X"FF",
  X"BF",  X"60",  X"60",  X"60",  X"40",  X"60",  X"BF",  X"05",
  X"BF",  X"20",  X"BF",  X"40",  X"FE",  X"BF",  X"BF",  X"00",
  X"06",  X"00",  X"BF",  X"20",  X"FE",  X"BF",  X"00",  X"00",
  X"20",  X"08",  X"20",  X"FF",  X"00",  X"E0",  X"BF",  X"BF",
  X"FE",  X"BF",  X"BF",  X"00",  X"20",  X"08",  X"20",  X"BF",
  X"BF",  X"FE",  X"BF",  X"A0",  X"20",  X"FD",  X"80",  X"20",
  X"20",  X"BF",  X"FD",  X"20",  X"BF",  X"00",  X"BF",  X"BF",
  X"08",  X"00",  X"BF",  X"00",  X"FD",  X"BF",  X"FE",  X"E0",
  X"A0",  X"FD",  X"00",  X"20",  X"20",  X"08",  X"00",  X"00",
  X"00",  X"05",  X"00",  X"20",  X"FF",  X"BF",  X"FD",  X"00",
  X"BF",  X"BF",  X"08",  X"00",  X"BF",  X"00",  X"FD",  X"BF",
  X"BF",  X"20",  X"00",  X"BF",  X"64",  X"BF",  X"FE",  X"BF",
  X"A0",  X"00",  X"00",  X"20",  X"07",  X"00",  X"00",  X"05",
  X"00",  X"20",  X"00",  X"BF",  X"A0",  X"00",  X"A0",  X"BF",
  X"BF",  X"80",  X"FE",  X"A0",  X"00",  X"BF",  X"BF",  X"60",
  X"FE",  X"BF",  X"00",  X"60",  X"00",  X"BF",  X"60",  X"FF",
  X"BF",  X"FE",  X"00",  X"A0",  X"FE",  X"40",  X"E0",  X"BF",
  X"BF",  X"06",  X"00",  X"BF",  X"A0",  X"A0",  X"00",  X"A0",
  X"20",  X"04",  X"A0",  X"00",  X"00",  X"07",  X"20",  X"BF",
  X"FD",  X"00",  X"20",  X"BF",  X"80",  X"FE",  X"BF",  X"BF",
  X"20",  X"00",  X"BF",  X"20",  X"80",  X"FE",  X"A0",  X"20",
  X"80",  X"FE",  X"A0",  X"20",  X"FF",  X"BF",  X"20",  X"40",
  X"60",  X"00",  X"80",  X"FE",  X"A0",  X"FF",  X"BF",  X"BF",
  X"60",  X"FF",  X"80",  X"FF",  X"BF",  X"A0",  X"20",  X"20",
  X"FC",  X"40",  X"FD",  X"60",  X"FD",  X"60",  X"BF",  X"20",
  X"00",  X"00",  X"20",  X"62",  X"00",  X"00",  X"00",  X"62",
  X"20",  X"00",  X"20",  X"20",  X"60",  X"00",  X"00",  X"20",
  X"E0",  X"60",  X"A0",  X"00",  X"60",  X"20",  X"60",  X"00",
  X"A0",  X"00",  X"00",  X"00",  X"00",  X"20",  X"20",  X"20",
  X"00",  X"20",  X"00",  X"E2",  X"00",  X"20",  X"00",  X"20",
  X"20",  X"20",  X"00",  X"40",  X"00",  X"20",  X"FF",  X"40",
  X"20",  X"A0",  X"3F",  X"A2",  X"00",  X"20",  X"0F",  X"20",
  X"00",  X"3F",  X"60",  X"62",  X"00",  X"20",  X"E0",  X"00",
  X"E2",  X"FF",  X"20",  X"0F",  X"20",  X"20",  X"E0",  X"00",
  X"0F",  X"20",  X"FF",  X"00",  X"00",  X"00",  X"FF",  X"20",
  X"60",  X"00",  X"02",  X"60",  X"00",  X"00",  X"63",  X"C0",
  X"02",  X"40",  X"00",  X"00",  X"60",  X"C0",  X"FF",  X"40",
  X"00",  X"BF",  X"20",  X"62",  X"00",  X"00",  X"0F",  X"20",
  X"E0",  X"20",  X"00",  X"20",  X"C0",  X"0F",  X"40",  X"00",
  X"BF",  X"00",  X"62",  X"00",  X"02",  X"61",  X"FF",  X"00",
  X"00",  X"BF",  X"20",  X"62",  X"00",  X"00",  X"0F",  X"20",
  X"E0",  X"20",  X"00",  X"20",  X"C0",  X"0F",  X"40",  X"00",
  X"BF",  X"FF",  X"00",  X"00",  X"62",  X"02",  X"62",  X"00",
  X"BF",  X"00",  X"62",  X"20",  X"00",  X"62",  X"20",  X"00",
  X"62",  X"20",  X"20",  X"20",  X"20",  X"00",  X"20",  X"20",
  X"20",  X"20",  X"20",  X"00",  X"62",  X"20",  X"BF",  X"0F",
  X"00",  X"00",  X"0F",  X"20",  X"00",  X"0F",  X"20",  X"0F",
  X"00",  X"E0",  X"00",  X"BF",  X"00",  X"61",  X"20",  X"20",
  X"20",  X"20",  X"20",  X"22",  X"22",  X"22",  X"22",  X"00",
  X"20",  X"FF",  X"20",  X"20",  X"00",  X"00",  X"20",  X"FF",
  X"20",  X"20",  X"20",  X"FF",  X"20",  X"00",  X"BF",  X"60",
  X"60",  X"00",  X"20",  X"00",  X"00",  X"EE",  X"20",  X"20",
  X"00",  X"20",  X"20",  X"00",  X"20",  X"00",  X"03",  X"20",
  X"E0",  X"00",  X"BF",  X"FF",  X"00",  X"00",  X"60",  X"60",
  X"60",  X"00",  X"00",  X"62",  X"60",  X"7F",  X"00",  X"60",
  X"00",  X"40",  X"00",  X"20",  X"20",  X"A0",  X"FF",  X"7F",
  X"3F",  X"20",  X"20",  X"20",  X"BF",  X"0F",  X"00",  X"20",
  X"0F",  X"00",  X"00",  X"0E",  X"20",  X"0F",  X"00",  X"FF",
  X"00",  X"00",  X"20",  X"20",  X"20",  X"20",  X"20",  X"20",
  X"20",  X"20",  X"20",  X"E0",  X"00",  X"40",  X"20",  X"00",
  X"00",  X"FF",  X"00",  X"FF",  X"00",  X"FF",  X"62",  X"FF",
  X"20",  X"20",  X"FF",  X"40",  X"FF",  X"20",  X"20",  X"FF",
  X"00",  X"BF",  X"EF",  X"00",  X"00",  X"20",  X"20",  X"60",
  X"7F",  X"6F",  X"40",  X"70",  X"70",  X"6F",  X"00",  X"00",
  X"EF",  X"20",  X"20",  X"40",  X"00",  X"00",  X"00",  X"00",
  X"EF",  X"20",  X"E0",  X"00",  X"EF",  X"00",  X"3F",  X"00",
  X"40",  X"20",  X"60",  X"00",  X"A0",  X"00",  X"20",  X"62",
  X"80",  X"EF",  X"62",  X"E0",  X"00",  X"00",  X"EF",  X"20",
  X"20",  X"00",  X"A0",  X"FF",  X"00",  X"E0",  X"00",  X"00",
  X"A0",  X"E2",  X"FF",  X"60",  X"BF",  X"60",  X"00",  X"00",
  X"EF",  X"00",  X"7F",  X"A0",  X"3F",  X"00",  X"80",  X"20",
  X"E0",  X"20",  X"C0",  X"00",  X"7F",  X"E0",  X"20",  X"00",
  X"20",  X"7F",  X"80",  X"40",  X"A0",  X"20",  X"C0",  X"00",
  X"20",  X"A0",  X"E0",  X"20",  X"A0",  X"C0",  X"E0",  X"E0",
  X"00",  X"60",  X"20",  X"00",  X"40",  X"E0",  X"E0",  X"60",
  X"E0",  X"60",  X"80",  X"20",  X"00",  X"A0",  X"61",  X"00",
  X"60",  X"60",  X"E0",  X"00",  X"E0",  X"60",  X"20",  X"20",
  X"00",  X"60",  X"C0",  X"00",  X"E0",  X"00",  X"20",  X"40",
  X"00",  X"E0",  X"E0",  X"3F",  X"40",  X"FF",  X"E0",  X"E0",
  X"A0",  X"A0",  X"E0",  X"60",  X"EF",  X"00",  X"E0",  X"00",
  X"E0",  X"00",  X"E0",  X"40",  X"FF",  X"E0",  X"60",  X"60",
  X"80",  X"A0",  X"60",  X"A0",  X"A0",  X"EF",  X"00",  X"60",
  X"00",  X"E0",  X"A0",  X"A0",  X"20",  X"60",  X"E0",  X"60",
  X"20",  X"80",  X"00",  X"20",  X"EF",  X"00",  X"20",  X"00",
  X"40",  X"7F",  X"80",  X"A0",  X"A0",  X"40",  X"60",  X"E0",
  X"20",  X"60",  X"A0",  X"00",  X"A0",  X"40",  X"FF",  X"00",
  X"62",  X"FF",  X"00",  X"EF",  X"00",  X"E0",  X"FF",  X"20",
  X"E0",  X"00",  X"E1",  X"60",  X"20",  X"FF",  X"20",  X"20",
  X"20",  X"40",  X"40",  X"20",  X"FF",  X"00",  X"00",  X"E5",
  X"60",  X"20",  X"FF",  X"20",  X"23",  X"FF",  X"20",  X"60",
  X"20",  X"FF",  X"20",  X"BF",  X"60",  X"60",  X"00",  X"00",
  X"20",  X"A0",  X"00",  X"00",  X"20",  X"E0",  X"00",  X"00",
  X"A0",  X"40",  X"20",  X"00",  X"20",  X"A0",  X"00",  X"00",
  X"A4",  X"00",  X"00",  X"24",  X"20",  X"40",  X"20",  X"20",
  X"00",  X"80",  X"60",  X"40",  X"60",  X"00",  X"60",  X"C0",
  X"A0",  X"FF",  X"00",  X"40",  X"60",  X"FF",  X"60",  X"20",
  X"E0",  X"00",  X"00",  X"A0",  X"A2",  X"00",  X"20",  X"20",
  X"20",  X"20",  X"E0",  X"00",  X"40",  X"E0",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"20",  X"20",  X"80",  X"40",
  X"00",  X"00",  X"20",  X"00",  X"00",  X"40",  X"00",  X"02",
  X"00",  X"00",  X"40",  X"00",  X"FD",  X"00",  X"20",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"60",  X"40",  X"60",  X"FF",
  X"60",  X"C0",  X"E0",  X"FF",  X"80",  X"40",  X"60",  X"20",
  X"FF",  X"60",  X"00",  X"80",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"02",  X"00",  X"20",  X"00",  X"80",  X"40",  X"20",
  X"00",  X"00",  X"00",  X"60",  X"40",  X"E0",  X"FF",  X"60",
  X"20",  X"80",  X"00",  X"A0",  X"00",  X"40",  X"60",  X"60",
  X"62",  X"00",  X"20",  X"80",  X"FF",  X"00",  X"60",  X"FF",
  X"00",  X"20",  X"00",  X"80",  X"40",  X"80",  X"06",  X"00",
  X"20",  X"00",  X"40",  X"20",  X"20",  X"00",  X"20",  X"00",
  X"FF",  X"00",  X"60",  X"FF",  X"60",  X"C0",  X"00",  X"00",
  X"00",  X"20",  X"00",  X"00",  X"20",  X"00",  X"01",  X"00",
  X"00",  X"40",  X"00",  X"FD",  X"00",  X"20",  X"FF",  X"60",
  X"20",  X"60",  X"20",  X"E0",  X"3F",  X"20",  X"80",  X"00",
  X"00",  X"20",  X"20",  X"40",  X"00",  X"20",  X"FF",  X"20",
  X"FF",  X"00",  X"01",  X"00",  X"20",  X"00",  X"80",  X"40",
  X"20",  X"00",  X"00",  X"FF",  X"00",  X"40",  X"00",  X"00",
  X"20",  X"20",  X"40",  X"00",  X"20",  X"FF",  X"20",  X"00",
  X"FF",  X"60",  X"FD",  X"00",  X"20",  X"FF",  X"20",  X"FF",
  X"60",  X"01",  X"00",  X"20",  X"00",  X"80",  X"40",  X"20",
  X"00",  X"FF",  X"00",  X"20",  X"00",  X"01",  X"E0",  X"20",
  X"FF",  X"20",  X"20",  X"FF",  X"00",  X"00",  X"F7",  X"3F",
  X"20",  X"FF",  X"00",  X"20",  X"FF",  X"00",  X"80",  X"FE",
  X"20",  X"FF",  X"20",  X"BF",  X"FD",  X"00",  X"22",  X"00",
  X"20",  X"E0",  X"BF",  X"00",  X"E0",  X"00",  X"C0",  X"60",
  X"00",  X"BF",  X"00",  X"00",  X"40",  X"00",  X"60",  X"00",
  X"62",  X"00",  X"60",  X"BF",  X"00",  X"C0",  X"60",  X"60",
  X"60",  X"A0",  X"FF",  X"BF",  X"A0",  X"A2",  X"FF",  X"60",
  X"60",  X"0C",  X"00",  X"60",  X"60",  X"FF",  X"60",  X"0C",
  X"00",  X"BF",  X"FF",  X"60",  X"C0",  X"E0",  X"FF",  X"E0",
  X"FD",  X"00",  X"E0",  X"00",  X"BF",  X"FD",  X"00",  X"22",
  X"00",  X"20",  X"A0",  X"7F",  X"00",  X"A0",  X"00",  X"80",
  X"20",  X"BF",  X"00",  X"00",  X"40",  X"00",  X"20",  X"00",
  X"62",  X"00",  X"20",  X"7F",  X"00",  X"80",  X"20",  X"20",
  X"60",  X"A0",  X"FF",  X"7F",  X"A0",  X"A2",  X"FF",  X"20",
  X"20",  X"0C",  X"00",  X"20",  X"60",  X"FF",  X"20",  X"0C",
  X"00",  X"7F",  X"FF",  X"20",  X"80",  X"A0",  X"FF",  X"A0",
  X"FC",  X"00",  X"E0",  X"00",  X"00",  X"E0",  X"61",  X"00",
  X"E0",  X"21",  X"00",  X"E0",  X"21",  X"BF",  X"00",  X"A0",
  X"00",  X"00",  X"20",  X"00",  X"00",  X"07",  X"00",  X"20",
  X"00",  X"00",  X"20",  X"20",  X"E0",  X"60",  X"00",  X"20",
  X"07",  X"60",  X"20",  X"FF",  X"20",  X"E0",  X"00",  X"00",
  X"00",  X"A2",  X"00",  X"00",  X"C0",  X"FF",  X"40",  X"00",
  X"BF",  X"20",  X"60",  X"00",  X"20",  X"20",  X"60",  X"00",
  X"00",  X"22",  X"08",  X"BF",  X"20",  X"00",  X"BF",  X"00",
  X"80",  X"00",  X"40",  X"00",  X"00",  X"3F",  X"40",  X"00",
  X"20",  X"20",  X"68",  X"00",  X"20",  X"20",  X"68",  X"20",
  X"20",  X"22",  X"EB",  X"24",  X"20",  X"00",  X"00",  X"20",
  X"62",  X"A0",  X"20",  X"00",  X"20",  X"00",  X"A1",  X"60",
  X"24",  X"60",  X"00",  X"20",  X"09",  X"20",  X"20",  X"00",
  X"00",  X"20",  X"60",  X"20",  X"E0",  X"00",  X"20",  X"00",
  X"20",  X"20",  X"E0",  X"00",  X"00",  X"62",  X"80",  X"FF",
  X"20",  X"64",  X"24",  X"20",  X"FF",  X"20",  X"20",  X"A0",
  X"20",  X"20",  X"00",  X"20",  X"20",  X"20",  X"E0",  X"00",
  X"BF",  X"60",  X"A0",  X"00",  X"00",  X"20",  X"00",  X"60",
  X"BF",  X"40",  X"20",  X"60",  X"22",  X"40",  X"E0",  X"60",
  X"40",  X"00",  X"40",  X"40",  X"80",  X"40",  X"00",  X"BF",
  X"00",  X"40",  X"00",  X"00",  X"20",  X"40",  X"00",  X"20",
  X"20",  X"40",  X"00",  X"20",  X"20",  X"40",  X"00",  X"20",
  X"A0",  X"FF",  X"20",  X"00",  X"A0",  X"00",  X"40",  X"E0",
  X"20",  X"A0",  X"FF",  X"60",  X"40",  X"80",  X"FF",  X"BF",
  X"E0",  X"00",  X"E0",  X"00",  X"BF",  X"A0",  X"00",  X"00",
  X"00",  X"00",  X"40",  X"60",  X"00",  X"00",  X"E0",  X"00",
  X"20",  X"00",  X"40",  X"60",  X"40",  X"FF",  X"00",  X"E0",
  X"00",  X"00",  X"80",  X"40",  X"FF",  X"E0",  X"A0",  X"60",
  X"A0",  X"60",  X"A0",  X"60",  X"A0",  X"FF",  X"60",  X"BF",
  X"A0",  X"60",  X"60",  X"80",  X"60",  X"A0",  X"40",  X"00",
  X"FF",  X"00",  X"20",  X"00",  X"40",  X"60",  X"80",  X"A0",
  X"FF",  X"00",  X"BF",  X"A0",  X"60",  X"60",  X"80",  X"60",
  X"00",  X"FF",  X"40",  X"BF",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"40",  X"00",  X"00",  X"A0",  X"A0",  X"00",  X"BF",
  X"00",  X"7F",  X"40",  X"BF",  X"FF",  X"FF",  X"FF",  X"80",
  X"E0",  X"00",  X"A0",  X"00",  X"40",  X"E0",  X"FF",  X"20",
  X"00",  X"40",  X"60",  X"40",  X"FF",  X"00",  X"E0",  X"00",
  X"60",  X"FF",  X"E0",  X"00",  X"00",  X"00",  X"80",  X"40",
  X"FF",  X"E0",  X"A0",  X"60",  X"A0",  X"60",  X"A0",  X"60",
  X"A0",  X"FF",  X"60",  X"BF",  X"A0",  X"60",  X"60",  X"80",
  X"60",  X"A0",  X"40",  X"00",  X"FF",  X"00",  X"20",  X"00",
  X"40",  X"60",  X"80",  X"A0",  X"FF",  X"00",  X"BF",  X"A0",
  X"60",  X"60",  X"80",  X"60",  X"00",  X"FF",  X"40",  X"BF",
  X"60",  X"A0",  X"00",  X"00",  X"20",  X"00",  X"20",  X"E0",
  X"40",  X"A0",  X"60",  X"00",  X"80",  X"00",  X"00",  X"00",
  X"40",  X"60",  X"60",  X"60",  X"3F",  X"20",  X"FF",  X"60",
  X"BF",  X"60",  X"7F",  X"A0",  X"60",  X"00",  X"00",  X"20",
  X"40",  X"60",  X"80",  X"20",  X"FF",  X"40",  X"BF",  X"60",
  X"7F",  X"60",  X"40",  X"00",  X"A0",  X"00",  X"20",  X"80",
  X"60",  X"40",  X"FF",  X"80",  X"E0",  X"00",  X"60",  X"00",
  X"00",  X"20",  X"60",  X"60",  X"80",  X"40",  X"80",  X"E0",
  X"00",  X"00",  X"FF",  X"00",  X"00",  X"20",  X"60",  X"20",
  X"C0",  X"40",  X"00",  X"00",  X"20",  X"60",  X"40",  X"00",
  X"00",  X"20",  X"60",  X"40",  X"00",  X"60",  X"20",  X"60",
  X"60",  X"00",  X"00",  X"40",  X"00",  X"20",  X"E0",  X"00",
  X"E0",  X"20",  X"00",  X"60",  X"00",  X"00",  X"60",  X"00",
  X"20",  X"60",  X"00",  X"20",  X"60",  X"00",  X"E0",  X"00",
  X"A3",  X"40",  X"00",  X"20",  X"60",  X"00",  X"60",  X"A0",
  X"60",  X"60",  X"00",  X"60",  X"A0",  X"60",  X"60",  X"00",
  X"60",  X"A0",  X"60",  X"60",  X"00",  X"00",  X"60",  X"60",
  X"00",  X"A0",  X"00",  X"E0",  X"00",  X"60",  X"60",  X"FF",
  X"20",  X"FF",  X"A0",  X"20",  X"E0",  X"00",  X"60",  X"20",
  X"00",  X"E0",  X"00",  X"BF",  X"00",  X"60",  X"20",  X"00",
  X"00",  X"A0",  X"A0",  X"40",  X"40",  X"E0",  X"A0",  X"60",
  X"BF",  X"FF",  X"80",  X"C0",  X"40",  X"00",  X"40",  X"FF",
  X"BF",  X"E0",  X"00",  X"40",  X"20",  X"20",  X"E0",  X"00",
  X"FC",  X"30",  X"00",  X"40",  X"60",  X"00",  X"BF",  X"00",
  X"20",  X"A0",  X"A0",  X"E0",  X"BF",  X"00",  X"60",  X"60",
  X"00",  X"02",  X"7F",  X"60",  X"00",  X"20",  X"20",  X"00",
  X"A0",  X"A0",  X"E0",  X"BF",  X"00",  X"20",  X"00",  X"FF",
  X"00",  X"20",  X"00",  X"A0",  X"A0",  X"E0",  X"BF",  X"BF",
  X"20",  X"20",  X"20",  X"00",  X"FF",  X"00",  X"20",  X"40",
  X"40",  X"00",  X"20",  X"00",  X"20",  X"20",  X"00",  X"80",
  X"00",  X"20",  X"3F",  X"40",  X"40",  X"20",  X"FC",  X"40",
  X"40",  X"40",  X"BF",  X"BF",  X"E0",  X"00",  X"00",  X"00",
  X"20",  X"3F",  X"00",  X"FC",  X"20",  X"00",  X"80",  X"00",
  X"20",  X"3F",  X"00",  X"40",  X"40",  X"FC",  X"40",  X"00",
  X"00",  X"00",  X"BF",  X"BF",  X"E0",  X"00",  X"FC",  X"00",
  X"40",  X"BF",  X"BF",  X"E0",  X"00",  X"3F",  X"3F",  X"FF",
  X"3F",  X"FF",  X"20",  X"BF",  X"BF",  X"FF",  X"00",  X"00",
  X"BF",  X"00",  X"BF",  X"FF",  X"BF",  X"20",  X"60",  X"BF",
  X"BF",  X"00",  X"C0",  X"BF",  X"A0",  X"BF",  X"40",  X"60",
  X"00",  X"00",  X"BF",  X"60",  X"BF",  X"40",  X"BF",  X"BF",
  X"00",  X"09",  X"E0",  X"00",  X"BF",  X"60",  X"BF",  X"80",
  X"BF",  X"BF",  X"00",  X"09",  X"E0",  X"00",  X"20",  X"00",
  X"00",  X"61",  X"00",  X"61",  X"3F",  X"FF",  X"09",  X"E0",
  X"00",  X"20",  X"00",  X"61",  X"E0",  X"40",  X"BF",  X"20",
  X"60",  X"00",  X"00",  X"60",  X"40",  X"20",  X"00",  X"00",
  X"00",  X"40",  X"20",  X"20",  X"E0",  X"00",  X"00",  X"20",
  X"04",  X"20",  X"20",  X"00",  X"20",  X"FF",  X"20",  X"E0",
  X"00",  X"20",  X"20",  X"00",  X"20",  X"04",  X"A0",  X"20",
  X"FF",  X"00",  X"20",  X"20",  X"20",  X"20",  X"E0",  X"00",
  X"BF",  X"20",  X"00",  X"BF",  X"FF",  X"BF",  X"FC",  X"40",
  X"BF",  X"00",  X"00",  X"40",  X"60",  X"A0",  X"00",  X"00",
  X"04",  X"80",  X"BF",  X"60",  X"00",  X"00",  X"BF",  X"FE",
  X"BF",  X"20",  X"00",  X"BF",  X"BF",  X"20",  X"BF",  X"00",
  X"20",  X"20",  X"20",  X"A0",  X"00",  X"20",  X"3B",  X"20",
  X"C0",  X"60",  X"00",  X"FE",  X"60",  X"20",  X"00",  X"00",
  X"E0",  X"00",  X"FE",  X"BF",  X"BF",  X"20",  X"20",  X"20",
  X"20",  X"A0",  X"FF",  X"20",  X"BB",  X"80",  X"C0",  X"20",
  X"40",  X"00",  X"E0",  X"00",  X"BF",  X"00",  X"40",  X"80",
  X"20",  X"40",  X"FF",  X"BF",  X"BF",  X"60",  X"A0",  X"40",
  X"00",  X"00",  X"60",  X"00",  X"00",  X"20",  X"60",  X"FF",
  X"60",  X"60",  X"A0",  X"20",  X"20",  X"60",  X"60",  X"40",
  X"60",  X"00",  X"80",  X"60",  X"60",  X"23",  X"A0",  X"20",
  X"20",  X"80",  X"00",  X"60",  X"40",  X"E0",  X"C0",  X"80",
  X"C0",  X"C0",  X"E0",  X"C0",  X"60",  X"A0",  X"40",  X"20",
  X"60",  X"40",  X"FF",  X"A0",  X"00",  X"00",  X"7F",  X"00",
  X"23",  X"00",  X"E0",  X"C0",  X"80",  X"E0",  X"80",  X"60",
  X"20",  X"40",  X"40",  X"60",  X"FF",  X"A0",  X"7F",  X"A0",
  X"00",  X"7F",  X"7F",  X"40",  X"A0",  X"FF",  X"3F",  X"20",
  X"E0",  X"00",  X"60",  X"60",  X"60",  X"80",  X"40",  X"A0",
  X"60",  X"7F",  X"BF",  X"40",  X"80",  X"00",  X"00",  X"00",
  X"FF",  X"7F",  X"FF",  X"20",  X"20",  X"20",  X"20",  X"E0",
  X"00",  X"00",  X"FF",  X"00",  X"20",  X"00",  X"00",  X"FF",
  X"60",  X"BF",  X"60",  X"60",  X"20",  X"A0",  X"00",  X"00",
  X"00",  X"00",  X"60",  X"60",  X"00",  X"FF",  X"60",  X"FF",
  X"00",  X"60",  X"00",  X"20",  X"20",  X"40",  X"A0",  X"80",
  X"FF",  X"60",  X"A0",  X"60",  X"00",  X"60",  X"60",  X"20",
  X"A0",  X"20",  X"60",  X"40",  X"00",  X"20",  X"20",  X"20",
  X"00",  X"80",  X"40",  X"C0",  X"40",  X"60",  X"80",  X"A0",
  X"00",  X"FF",  X"C0",  X"40",  X"00",  X"00",  X"A0",  X"60",
  X"60",  X"80",  X"40",  X"3F",  X"80",  X"20",  X"E0",  X"00",
  X"80",  X"40",  X"A0",  X"00",  X"FF",  X"60",  X"80",  X"40",
  X"A0",  X"00",  X"FF",  X"60",  X"FF",  X"A0",  X"BF",  X"60",
  X"A0",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"60",
  X"00",  X"80",  X"00",  X"60",  X"60",  X"FE",  X"A0",  X"20",
  X"E0",  X"00",  X"E0",  X"C0",  X"00",  X"00",  X"00",  X"40",
  X"60",  X"C0",  X"FF",  X"40",  X"60",  X"60",  X"40",  X"60",
  X"BF",  X"20",  X"A0",  X"20",  X"80",  X"20",  X"40",  X"00",
  X"60",  X"00",  X"63",  X"40",  X"40",  X"00",  X"BF",  X"BF",
  X"00",  X"20",  X"80",  X"BF",  X"04",  X"00",  X"00",  X"BF",
  X"C0",  X"00",  X"04",  X"20",  X"80",  X"E0",  X"A0",  X"00",
  X"C0",  X"20",  X"A0",  X"00",  X"40",  X"20",  X"FF",  X"60",
  X"00",  X"40",  X"60",  X"60",  X"00",  X"BF",  X"C0",  X"BF",
  X"00",  X"00",  X"20",  X"80",  X"BF",  X"00",  X"04",  X"A0",
  X"C0",  X"C0",  X"20",  X"BF",  X"00",  X"20",  X"04",  X"E0",
  X"20",  X"00",  X"A0",  X"80",  X"40",  X"00",  X"40",  X"FF",
  X"60",  X"00",  X"60",  X"00",  X"FF",  X"E0",  X"A0",  X"00",
  X"20",  X"FF",  X"60",  X"00",  X"FF",  X"20",  X"E0",  X"00",
  X"C0",  X"60",  X"00",  X"20",  X"BF",  X"FF",  X"FF",  X"20",
  X"E0",  X"00",  X"00",  X"00",  X"FF",  X"00",  X"BF",  X"20",
  X"FE",  X"00",  X"20",  X"20",  X"20",  X"E0",  X"00",  X"BF",
  X"60",  X"00",  X"60",  X"63",  X"20",  X"40",  X"00",  X"03",
  X"00",  X"20",  X"C0",  X"03",  X"00",  X"E0",  X"C0",  X"C0",
  X"E0",  X"40",  X"40",  X"A0",  X"60",  X"00",  X"FF",  X"E0",
  X"E0",  X"00",  X"00",  X"60",  X"00",  X"00",  X"60",  X"20",
  X"60",  X"40",  X"20",  X"60",  X"60",  X"E0",  X"00",  X"60",
  X"FE",  X"00",  X"60",  X"00",  X"60",  X"A0",  X"20",  X"FC",
  X"A0",  X"20",  X"60",  X"60",  X"80",  X"40",  X"80",  X"FF",
  X"00",  X"BF",  X"A0",  X"00",  X"00",  X"A0",  X"A0",  X"00",
  X"00",  X"20",  X"60",  X"00",  X"00",  X"A0",  X"00",  X"00",
  X"A0",  X"A0",  X"00",  X"00",  X"40",  X"20",  X"00",  X"00",
  X"00",  X"A0",  X"FF",  X"A0",  X"00",  X"00",  X"FF",  X"00",
  X"60",  X"00",  X"A0",  X"20",  X"60",  X"60",  X"80",  X"40",
  X"80",  X"A0",  X"FF",  X"00",  X"E0",  X"00",  X"00",  X"FF",
  X"00",  X"40",  X"00",  X"FF",  X"00",  X"7F",  X"00",  X"60",
  X"A2",  X"80",  X"00",  X"00",  X"FF",  X"20",  X"FF",  X"00",
  X"FF",  X"22",  X"20",  X"00",  X"FF",  X"00",  X"BF",  X"20",
  X"03",  X"E0",  X"00",  X"20",  X"20",  X"00",  X"20",  X"60",
  X"00",  X"FF",  X"60",  X"FD",  X"00",  X"20",  X"20",  X"20",
  X"A0",  X"60",  X"00",  X"20",  X"60",  X"40",  X"00",  X"FF",
  X"00",  X"FF",  X"20",  X"60",  X"80",  X"FF",  X"40",  X"80",
  X"00",  X"BF",  X"C0",  X"00",  X"20",  X"80",  X"00",  X"FF",
  X"00",  X"FF",  X"20",  X"A0",  X"80",  X"C0",  X"FF",  X"80",
  X"E0",  X"00",  X"BF",  X"60",  X"00",  X"00",  X"E6",  X"00",
  X"E8",  X"00",  X"7F",  X"A0",  X"A0",  X"60",  X"00",  X"00",
  X"20",  X"20",  X"40",  X"00",  X"20",  X"E0",  X"20",  X"7F",
  X"00",  X"40",  X"FF",  X"60",  X"20",  X"FF",  X"BF",  X"C0",
  X"00",  X"00",  X"00",  X"20",  X"20",  X"80",  X"00",  X"00",
  X"60",  X"60",  X"7F",  X"40",  X"60",  X"60",  X"00",  X"20",
  X"7F",  X"40",  X"80",  X"00",  X"60",  X"A0",  X"00",  X"60",
  X"7F",  X"80",  X"E0",  X"00",  X"BF",  X"40",  X"00",  X"80",
  X"40",  X"80",  X"00",  X"60",  X"00",  X"80",  X"00",  X"00",
  X"E0",  X"E0",  X"FF",  X"E0",  X"A0",  X"A0",  X"00",  X"60",
  X"A0",  X"00",  X"00",  X"00",  X"40",  X"E0",  X"A0",  X"E0",
  X"60",  X"E0",  X"00",  X"60",  X"60",  X"E0",  X"A0",  X"E0",
  X"60",  X"E0",  X"00",  X"60",  X"40",  X"E0",  X"E0",  X"60",
  X"E0",  X"60",  X"40",  X"C0",  X"00",  X"00",  X"60",  X"E0",
  X"60",  X"E0",  X"00",  X"E0",  X"00",  X"A0",  X"80",  X"E0",
  X"00",  X"80",  X"60",  X"40",  X"A0",  X"80",  X"A0",  X"60",
  X"A0",  X"E7",  X"00",  X"E0",  X"00",  X"60",  X"40",  X"A0",
  X"E0",  X"60",  X"40",  X"00",  X"60",  X"A0",  X"60",  X"F8",
  X"60",  X"FF",  X"FF",  X"20",  X"60",  X"A0",  X"00",  X"20",
  X"00",  X"FF",  X"E0",  X"80",  X"60",  X"40",  X"40",  X"FF",
  X"80",  X"E0",  X"E0",  X"FF",  X"E0",  X"A0",  X"A0",  X"00",
  X"60",  X"A0",  X"00",  X"00",  X"00",  X"40",  X"E0",  X"A0",
  X"E0",  X"60",  X"E0",  X"00",  X"60",  X"60",  X"E0",  X"A0",
  X"E0",  X"60",  X"E0",  X"00",  X"60",  X"40",  X"E0",  X"E0",
  X"60",  X"E0",  X"60",  X"40",  X"80",  X"60",  X"A0",  X"60",
  X"A0",  X"C0",  X"40",  X"A0",  X"60",  X"20",  X"00",  X"E0",
  X"60",  X"40",  X"E7",  X"E0",  X"E0",  X"00",  X"00",  X"E5",
  X"00",  X"20",  X"00",  X"3F",  X"A0",  X"7F",  X"80",  X"80",
  X"00",  X"FF",  X"A0",  X"00",  X"A0",  X"00",  X"00",  X"00",
  X"40",  X"00",  X"A0",  X"20",  X"60",  X"20",  X"00",  X"60",
  X"60",  X"20",  X"A0",  X"20",  X"60",  X"20",  X"00",  X"60",
  X"60",  X"20",  X"60",  X"20",  X"60",  X"20",  X"80",  X"40",
  X"A0",  X"60",  X"A0",  X"60",  X"00",  X"F7",  X"00",  X"E7",
  X"00",  X"E0",  X"00",  X"60",  X"FF",  X"E0",  X"A0",  X"60",
  X"A0",  X"E0",  X"E0",  X"A0",  X"FF",  X"60",  X"00",  X"FA",
  X"00",  X"00",  X"FF",  X"E0",  X"20",  X"7F",  X"40",  X"40",
  X"FF",  X"00",  X"80",  X"40",  X"A0",  X"60",  X"20",  X"00",
  X"A0",  X"60",  X"40",  X"E7",  X"A0",  X"E0",  X"00",  X"FA",
  X"00",  X"FF",  X"00",  X"FF",  X"80",  X"A0",  X"BF",  X"00",
  X"80",  X"FF",  X"A0",  X"00",  X"FA",  X"00",  X"FF",  X"C0",
  X"BF",  X"20",  X"00",  X"00",  X"21",  X"A0",  X"00",  X"20",
  X"A0",  X"7F",  X"00",  X"80",  X"60",  X"60",  X"80",  X"40",
  X"40",  X"7F",  X"3F",  X"FF",  X"40",  X"80",  X"A0",  X"FF",
  X"A0",  X"20",  X"60",  X"00",  X"00",  X"40",  X"00",  X"E0",
  X"00",  X"FF",  X"62",  X"BF",  X"40",  X"60",  X"00",  X"00",
  X"FF",  X"00",  X"F7",  X"00",  X"00",  X"BF",  X"00",  X"62",
  X"00",  X"00",  X"00",  X"20",  X"60",  X"00",  X"21",  X"20",
  X"40",  X"20",  X"00",  X"60",  X"00",  X"00",  X"F7",  X"00",
  X"20",  X"FF",  X"00",  X"20",  X"60",  X"60",  X"FF",  X"40",
  X"F7",  X"00",  X"21",  X"20",  X"00",  X"20",  X"21",  X"00",
  X"00",  X"20",  X"00",  X"00",  X"F7",  X"00",  X"40",  X"FF",
  X"00",  X"20",  X"60",  X"00",  X"20",  X"F7",  X"00",  X"20",
  X"60",  X"00",  X"20",  X"E0",  X"00",  X"40",  X"00",  X"22",
  X"60",  X"FF",  X"00",  X"FF",  X"00",  X"00",  X"00",  X"FC",
  X"40",  X"00",  X"60",  X"00",  X"40",  X"80",  X"00",  X"00",
  X"60",  X"E0",  X"20",  X"00",  X"00",  X"00",  X"00",  X"20",
  X"00",  X"FC",  X"40",  X"E0",  X"20",  X"20",  X"00",  X"62",
  X"C0",  X"00",  X"40",  X"00",  X"BF",  X"00",  X"20",  X"62",
  X"00",  X"01",  X"00",  X"3F",  X"00",  X"00",  X"20",  X"80",
  X"20",  X"20",  X"E0",  X"00",  X"20",  X"00",  X"40",  X"20",
  X"E0",  X"00",  X"BF",  X"20",  X"00",  X"61",  X"00",  X"00",
  X"00",  X"00",  X"A2",  X"20",  X"20",  X"01",  X"20",  X"20",
  X"00",  X"40",  X"A2",  X"20",  X"20",  X"00",  X"00",  X"00",
  X"BF",  X"00",  X"20",  X"62",  X"00",  X"01",  X"00",  X"20",
  X"00",  X"20",  X"20",  X"40",  X"20",  X"E0",  X"00",  X"00",
  X"40",  X"20",  X"E0",  X"00",  X"40",  X"60",  X"00",  X"00",
  X"00",  X"40",  X"40",  X"00",  X"BF",  X"20",  X"A2",  X"E0",
  X"00",  X"40",  X"80",  X"40",  X"00",  X"20",  X"E0",  X"20",
  X"80",  X"40",  X"00",  X"20",  X"20",  X"60",  X"00",  X"40",
  X"40",  X"FF",  X"40",  X"00",  X"60",  X"00",  X"00",  X"00",
  X"40",  X"20",  X"00",  X"60",  X"60",  X"00",  X"00",  X"40",
  X"40",  X"FF",  X"40",  X"E0",  X"60",  X"E0",  X"C0",  X"40",
  X"E0",  X"60",  X"E0",  X"C0",  X"E0",  X"00",  X"BF",  X"20",
  X"00",  X"00",  X"00",  X"BF",  X"62",  X"40",  X"80",  X"20",
  X"20",  X"40",  X"00",  X"00",  X"60",  X"40",  X"80",  X"C0",
  X"80",  X"00",  X"40",  X"60",  X"40",  X"80",  X"C0",  X"80",
  X"FF",  X"60",  X"00",  X"40",  X"40",  X"A0",  X"FF",  X"60",
  X"40",  X"E0",  X"00",  X"BF",  X"00",  X"00",  X"00",  X"21",
  X"02",  X"00",  X"3F",  X"00",  X"21",  X"E0",  X"00",  X"60",
  X"FF",  X"00",  X"00",  X"E0",  X"00",  X"BF",  X"00",  X"00",
  X"00",  X"00",  X"E4",  X"00",  X"20",  X"00",  X"00",  X"3F",
  X"BF",  X"BF",  X"A0",  X"00",  X"A0",  X"00",  X"00",  X"00",
  X"20",  X"A0",  X"00",  X"20",  X"20",  X"20",  X"A0",  X"00",
  X"20",  X"20",  X"20",  X"20",  X"60",  X"40",  X"60",  X"E0",
  X"00",  X"F9",  X"20",  X"E0",  X"00",  X"BF",  X"00",  X"00",
  X"02",  X"21",  X"3F",  X"00",  X"21",  X"E0",  X"00",  X"60",
  X"FF",  X"00",  X"00",  X"E0",  X"00",  X"BF",  X"60",  X"00",
  X"20",  X"F5",  X"60",  X"60",  X"62",  X"00",  X"00",  X"00",
  X"62",  X"20",  X"00",  X"60",  X"20",  X"60",  X"00",  X"00",
  X"60",  X"60",  X"60",  X"00",  X"60",  X"60",  X"00",  X"20",
  X"60",  X"60",  X"00",  X"60",  X"40",  X"60",  X"20",  X"00",
  X"3F",  X"60",  X"60",  X"00",  X"60",  X"60",  X"60",  X"00",
  X"60",  X"40",  X"00",  X"60",  X"F5",  X"62",  X"60",  X"60",
  X"60",  X"00",  X"60",  X"F5",  X"62",  X"60",  X"60",  X"04",
  X"00",  X"04",  X"00",  X"F4",  X"00",  X"E0",  X"00",  X"04",
  X"00",  X"FF",  X"00",  X"04",  X"00",  X"F4",  X"20",  X"E0",
  X"00",  X"F5",  X"00",  X"60",  X"60",  X"60",  X"FF",  X"60",
  X"FF",  X"F5",  X"00",  X"FF",  X"60",  X"F4",  X"00",  X"FF",
  X"00",  X"00",  X"00",  X"62",  X"C0",  X"FF",  X"40",  X"00",
  X"BF",  X"00",  X"00",  X"00",  X"01",  X"21",  X"3F",  X"00",
  X"21",  X"E0",  X"00",  X"60",  X"FF",  X"00",  X"00",  X"E0",
  X"00",  X"BF",  X"00",  X"00",  X"00",  X"21",  X"01",  X"00",
  X"3F",  X"00",  X"21",  X"E0",  X"00",  X"60",  X"FF",  X"00",
  X"00",  X"E0",  X"00",  X"BF",  X"00",  X"00",  X"00",  X"21",
  X"01",  X"00",  X"3F",  X"00",  X"21",  X"E0",  X"00",  X"60",
  X"FF",  X"00",  X"00",  X"E0",  X"00",  X"00",  X"00",  X"2F",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"E0",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"20",  X"60",  X"E0",  X"40",  X"00",
  X"20",  X"40",  X"00",  X"40",  X"40",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"40",  X"00",  X"00",  X"20",  X"E0",  X"00",
  X"C0",  X"00",  X"00",  X"00",  X"C0",  X"00",  X"00",  X"40",
  X"00",  X"20",  X"60",  X"FF",  X"20",  X"40",  X"00",  X"A0",
  X"60",  X"60",  X"40",  X"00",  X"A0",  X"40",  X"FF",  X"00",
  X"00",  X"00",  X"A0",  X"00",  X"00",  X"C0",  X"20",  X"00",
  X"00",  X"A0",  X"00",  X"60",  X"C0",  X"00",  X"A0",  X"C0",
  X"A0",  X"A0",  X"FF",  X"C0",  X"00",  X"60",  X"40",  X"FF",
  X"20",  X"00",  X"20",  X"C0",  X"A0",  X"00",  X"60",  X"C0",
  X"00",  X"60",  X"C0",  X"00",  X"60",  X"C0",  X"00",  X"60",
  X"C0",  X"00",  X"A0",  X"C0",  X"00",  X"A0",  X"C0",  X"00",
  X"60",  X"C0",  X"00",  X"A0",  X"C0",  X"00",  X"A0",  X"C0",
  X"00",  X"60",  X"C0",  X"00",  X"60",  X"C0",  X"00",  X"A0",
  X"C0",  X"00",  X"A0",  X"C0",  X"00",  X"60",  X"C0",  X"00",
  X"A0",  X"C0",  X"00",  X"A0",  X"C0",  X"00",  X"60",  X"C0",
  X"00",  X"60",  X"C0",  X"00",  X"60",  X"C0",  X"00",  X"BF",
  X"C0",  X"00",  X"BF",  X"C0",  X"00",  X"60",  X"C0",  X"00",
  X"BF",  X"C0",  X"00",  X"BF",  X"C0",  X"00",  X"60",  X"C0",
  X"00",  X"60",  X"C0",  X"00",  X"BF",  X"C0",  X"00",  X"BF",
  X"C0",  X"00",  X"60",  X"C0",  X"00",  X"BF",  X"C0",  X"00",
  X"BF",  X"20",  X"FF",  X"C0",  X"00",  X"A0",  X"C0",  X"00",
  X"00",  X"E0",  X"00",  X"00",  X"20",  X"40",  X"00",  X"00",
  X"40",  X"00",  X"00",  X"00",  X"00",  X"00",  X"40",  X"00",
  X"00",  X"20",  X"E0",  X"00",  X"C0",  X"00",  X"00",  X"00",
  X"C0",  X"00",  X"00",  X"40",  X"00",  X"20",  X"60",  X"FF",
  X"20",  X"40",  X"00",  X"A0",  X"60",  X"60",  X"40",  X"00",
  X"A0",  X"40",  X"FF",  X"00",  X"00",  X"00",  X"A0",  X"00",
  X"00",  X"C0",  X"20",  X"00",  X"00",  X"A0",  X"00",  X"60",
  X"C0",  X"00",  X"A0",  X"C0",  X"A0",  X"A0",  X"FF",  X"C0",
  X"00",  X"60",  X"40",  X"FF",  X"20",  X"00",  X"20",  X"C0",
  X"A0",  X"00",  X"60",  X"C0",  X"00",  X"60",  X"C0",  X"00",
  X"60",  X"C0",  X"00",  X"60",  X"C0",  X"00",  X"A0",  X"C0",
  X"00",  X"A0",  X"C0",  X"00",  X"60",  X"C0",  X"00",  X"A0",
  X"C0",  X"00",  X"A0",  X"C0",  X"00",  X"60",  X"C0",  X"00",
  X"60",  X"C0",  X"00",  X"A0",  X"C0",  X"00",  X"A0",  X"C0",
  X"00",  X"60",  X"C0",  X"00",  X"A0",  X"C0",  X"00",  X"A0",
  X"C0",  X"00",  X"60",  X"C0",  X"00",  X"60",  X"C0",  X"00",
  X"60",  X"C0",  X"00",  X"BF",  X"C0",  X"00",  X"BF",  X"C0",
  X"00",  X"60",  X"C0",  X"00",  X"BF",  X"C0",  X"00",  X"BF",
  X"C0",  X"00",  X"60",  X"C0",  X"00",  X"60",  X"C0",  X"00",
  X"BF",  X"C0",  X"00",  X"BF",  X"C0",  X"00",  X"60",  X"C0",
  X"00",  X"BF",  X"C0",  X"00",  X"BF",  X"20",  X"FF",  X"C0",
  X"00",  X"C0",  X"C0",  X"00",  X"00",  X"E0",  X"00",  X"E0",
  X"20",  X"00",  X"20",  X"60",  X"E0",  X"60",  X"E0",  X"20",
  X"BF",  X"04",  X"3F",  X"20",  X"00",  X"E0",  X"00",  X"BF",
  X"A0",  X"00",  X"20",  X"00",  X"00",  X"00",  X"20",  X"80",
  X"00",  X"00",  X"00",  X"00",  X"40",  X"20",  X"20",  X"20",
  X"FF",  X"20",  X"E0",  X"20",  X"E0",  X"00",  X"00",  X"A1",
  X"60",  X"00",  X"00",  X"40",  X"A1",  X"E0",  X"00",  X"61",
  X"40",  X"A1",  X"A1",  X"E0",  X"00",  X"BF",  X"A0",  X"00",
  X"20",  X"00",  X"40",  X"00",  X"20",  X"20",  X"80",  X"00",
  X"00",  X"40",  X"20",  X"20",  X"60",  X"FF",  X"00",  X"00",
  X"20",  X"40",  X"20",  X"00",  X"20",  X"20",  X"80",  X"FF",
  X"40",  X"E0",  X"00",  X"00",  X"62",  X"60",  X"C0",  X"A0",
  X"FF",  X"20",  X"40",  X"20",  X"00",  X"00",  X"E0",  X"00",
  X"C0",  X"A0",  X"FF",  X"20",  X"40",  X"E0",  X"00",  X"00",
  X"62",  X"E0",  X"E0",  X"00",  X"20",  X"80",  X"60",  X"FF",
  X"00",  X"C0",  X"E0",  X"00",  X"00",  X"00",  X"E0",  X"00",
  X"22",  X"C0",  X"00",  X"00",  X"40",  X"00",  X"00",  X"00",
  X"A0",  X"A0",  X"A0",  X"A0",  X"A0",  X"A0",  X"A0",  X"A0",
  X"00",  X"00",  X"40",  X"80",  X"00",  X"00",  X"00",  X"00",
  X"E0",  X"00",  X"62",  X"C0",  X"40",  X"40",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"A0",  X"A0",  X"A0",  X"A0",  X"A0",
  X"A0",  X"A0",  X"A0",  X"00",  X"00",  X"40",  X"80",  X"00",
  X"00",  X"23",  X"00",  X"00",  X"E1",  X"C0",  X"20",  X"00",
  X"00",  X"00",  X"BF",  X"BF",  X"BF",  X"BF",  X"BF",  X"BF",
  X"BF",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"E1",  X"C0",  X"A0",  X"60",  X"A0",  X"A0",  X"02",
  X"00",  X"00",  X"21",  X"20",  X"20",  X"20",  X"20",  X"20",
  X"20",  X"00",  X"00",  X"6F",  X"60",  X"00",  X"00",  X"00",
  X"00",  X"22",  X"00",  X"20",  X"20",  X"00",  X"00",  X"00",
  X"00",  X"FF",  X"00",  X"00",  X"22",  X"00",  X"20",  X"00",
  X"00",  X"00",  X"20",  X"00",  X"FF",  X"00",  X"00",  X"00",
  X"21",  X"20",  X"20",  X"20",  X"20",  X"20",  X"20",  X"20",
  X"00",  X"00",  X"00",  X"80",  X"A0",  X"2F",  X"00",  X"00",
  X"00",  X"00",  X"80",  X"A0",  X"60",  X"00",  X"2F",  X"00",
  X"20",  X"00",  X"60",  X"00",  X"2F",  X"2F",  X"40",  X"00",
  X"00",  X"60",  X"00",  X"00",  X"20",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"60",  X"00",  X"00",  X"20",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"60",  X"00",  X"00",  X"FF",  X"20",
  X"80",  X"A0",  X"20",  X"E0",  X"20",  X"20",  X"E0",  X"20",
  X"20",  X"E0",  X"20",  X"00",  X"00",  X"2F",  X"E0",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"C0",  X"00",  X"00",  X"20",
  X"00",  X"22",  X"00",  X"00",  X"62",  X"40",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"60",  X"60",  X"60",  X"60",
  X"60",  X"60",  X"60",  X"60",  X"60",  X"60",  X"60",  X"60",
  X"60",  X"60",  X"60",  X"60",  X"60",  X"00",  X"A2",  X"80",
  X"00",  X"00",  X"00",  X"20",  X"20",  X"20",  X"20",  X"20",
  X"20",  X"20",  X"20",  X"20",  X"20",  X"20",  X"20",  X"20",
  X"20",  X"20",  X"20",  X"20",  X"20",  X"00",  X"00",  X"00",
  X"40",  X"80",  X"E0",  X"00",  X"E0",  X"00",  X"E0",  X"00",
  X"A0",  X"00",  X"00",  X"A0",  X"00",  X"21",  X"00",  X"00",
  X"22",  X"00",  X"60",  X"00",  X"E0",  X"2F",  X"00",  X"00",
  X"22",  X"00",  X"00",  X"00",  X"6F",  X"60",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"A0",  X"2F",  X"60",  X"00",  X"00",
  X"00",  X"00",  X"22",  X"00",  X"60",  X"00",  X"02",  X"00",
  X"BF",  X"00",  X"60",  X"62",  X"60",  X"20",  X"00",  X"40",
  X"60",  X"00",  X"E0",  X"22",  X"00",  X"40",  X"C0",  X"00",
  X"00",  X"00",  X"40",  X"00",  X"40",  X"60",  X"60",  X"FF",
  X"80",  X"40",  X"40",  X"A0",  X"20",  X"E0",  X"00",  X"40",
  X"E0",  X"00",  X"20",  X"00",  X"62",  X"40",  X"60",  X"E0",
  X"40",  X"BF",  X"00",  X"A2",  X"60",  X"40",  X"00",  X"A2",
  X"20",  X"00",  X"00",  X"20",  X"00",  X"62",  X"40",  X"20",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"20",  X"A1",  X"61",
  X"00",  X"E0",  X"00",  X"A0",  X"80",  X"80",  X"A0",  X"00",
  X"20",  X"80",  X"00",  X"00",  X"20",  X"00",  X"40",  X"00",
  X"40",  X"60",  X"00",  X"80",  X"40",  X"00",  X"80",  X"7F",
  X"80",  X"20",  X"20",  X"00",  X"00",  X"00",  X"60",  X"FF",
  X"20",  X"00",  X"A0",  X"FF",  X"C0",  X"A0",  X"FF",  X"00",
  X"20",  X"20",  X"FF",  X"00",  X"E0",  X"00",  X"A0",  X"FF",
  X"20",  X"00",  X"00",  X"E0",  X"60",  X"60",  X"00",  X"00",
  X"62",  X"00",  X"20",  X"40",  X"00",  X"62",  X"00",  X"20",
  X"40",  X"00",  X"20",  X"20",  X"01",  X"00",  X"00",  X"00",
  X"00",  X"20",  X"FC",  X"40",  X"03",  X"40",  X"00",  X"20",
  X"20",  X"02",  X"00",  X"00",  X"00",  X"00",  X"02",  X"00",
  X"00",  X"62",  X"40",  X"00",  X"20",  X"20",  X"01",  X"00",
  X"00",  X"00",  X"00",  X"02",  X"00",  X"60",  X"00",  X"62",
  X"40",  X"00",  X"20",  X"20",  X"01",  X"00",  X"00",  X"00",
  X"00",  X"01",  X"00",  X"00",  X"62",  X"40",  X"60",  X"A0",
  X"A0",  X"60",  X"00",  X"E0",  X"00",  X"00",  X"62",  X"20",
  X"20",  X"E0",  X"00",  X"BF",  X"00",  X"61",  X"00",  X"60",
  X"00",  X"20",  X"00",  X"40",  X"00",  X"00",  X"E0",  X"00",
  X"BF",  X"00",  X"61",  X"60",  X"00",  X"20",  X"40",  X"00",
  X"00",  X"E0",  X"00",  X"BF",  X"00",  X"61",  X"60",  X"00",
  X"20",  X"40",  X"00",  X"00",  X"E0",  X"00",  X"BF",  X"00",
  X"61",  X"60",  X"00",  X"20",  X"40",  X"00",  X"00",  X"E0",
  X"00",  X"BF",  X"00",  X"61",  X"60",  X"00",  X"20",  X"40",
  X"00",  X"00",  X"E0",  X"00",  X"BF",  X"00",  X"61",  X"60",
  X"00",  X"20",  X"40",  X"00",  X"00",  X"E0",  X"00",  X"BF",
  X"00",  X"61",  X"60",  X"00",  X"20",  X"40",  X"00",  X"00",
  X"E0",  X"00",  X"BF",  X"00",  X"61",  X"00",  X"60",  X"00",
  X"20",  X"00",  X"40",  X"00",  X"00",  X"E0",  X"00",  X"00",
  X"00",  X"62",  X"40",  X"00",  X"00",  X"60",  X"40",  X"00",
  X"62",  X"40",  X"00",  X"00",  X"62",  X"40",  X"00",  X"00",
  X"60",  X"60",  X"60",  X"00",  X"00",  X"40",  X"60",  X"40",
  X"00",  X"00",  X"FF",  X"00",  X"DC",  X"00",  X"A0",  X"DC",
  X"00",  X"20",  X"20",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"20",  X"00",  X"00",  X"00",  X"00",  X"80",  X"A0",  X"E0",
  X"00",  X"E0",  X"00",  X"00",  X"E0",  X"60",  X"60",  X"00",
  X"00",  X"00",  X"22",  X"20",  X"00",  X"40",  X"00",  X"00",
  X"22",  X"20",  X"00",  X"00",  X"20",  X"E0",  X"60",  X"00",
  X"E2",  X"C0",  X"60",  X"00",  X"E2",  X"C0",  X"00",  X"E2",
  X"60",  X"C0",  X"E0",  X"00",  X"E0",  X"00",  X"20",  X"00",
  X"00",  X"00",  X"40",  X"80",  X"00",  X"60",  X"60",  X"60",
  X"00",  X"00",  X"40",  X"00",  X"40",  X"40",  X"00",  X"00",
  X"21",  X"00",  X"BF",  X"00",  X"00",  X"20",  X"60",  X"00",
  X"00",  X"00",  X"00",  X"20",  X"00",  X"20",  X"00",  X"00",
  X"00",  X"FF",  X"00",  X"E0",  X"00",  X"A1",  X"60",  X"60",
  X"60",  X"60",  X"60",  X"60",  X"60",  X"00",  X"60",  X"60",
  X"60",  X"60",  X"60",  X"00",  X"A2",  X"61",  X"60",  X"A2",
  X"20",  X"00",  X"00",  X"00",  X"00",  X"E0",  X"00",  X"E2",
  X"C0",  X"C0",  X"A0",  X"00",  X"A0",  X"A0",  X"A0",  X"A0",
  X"A0",  X"A0",  X"A0",  X"A0",  X"A0",  X"00",  X"A0",  X"00",
  X"00",  X"A1",  X"80",  X"80",  X"00",  X"00",  X"80",  X"A0",
  X"A1",  X"00",  X"E2",  X"20",  X"20",  X"40",  X"00",  X"A2",
  X"40",  X"40",  X"00",  X"80",  X"00",  X"A0",  X"00",  X"E2",
  X"80",  X"40",  X"60",  X"60",  X"A0",  X"60",  X"A0",  X"A0",
  X"A0",  X"A0",  X"A0",  X"A0",  X"A0",  X"A0",  X"A0",  X"A0",
  X"A0",  X"00",  X"A0",  X"A0",  X"A0",  X"A0",  X"A0",  X"A0",
  X"A0",  X"A0",  X"00",  X"00",  X"A0",  X"60",  X"A0",  X"A0",
  X"A0",  X"A0",  X"A0",  X"A0",  X"A0",  X"A0",  X"A0",  X"A0",
  X"A0",  X"20",  X"00",  X"00",  X"00",  X"40",  X"80",  X"A1",
  X"61",  X"00",  X"00",  X"60",  X"60",  X"60",  X"60",  X"00",
  X"60",  X"00",  X"A2",  X"61",  X"60",  X"A2",  X"E0",  X"20",
  X"00",  X"00",  X"00",  X"00",  X"E0",  X"00",  X"E2",  X"C0",
  X"C0",  X"A0",  X"00",  X"A0",  X"A0",  X"A0",  X"A0",  X"A0",
  X"A0",  X"A0",  X"A0",  X"A0",  X"00",  X"A0",  X"00",  X"00",
  X"A1",  X"80",  X"80",  X"00",  X"00",  X"80",  X"A0",  X"A1",
  X"00",  X"E2",  X"00",  X"E2",  X"80",  X"00",  X"00",  X"A1",
  X"00",  X"80",  X"00",  X"00",  X"00",  X"A0",  X"80",  X"00",
  X"00",  X"E2",  X"20",  X"20",  X"40",  X"00",  X"A2",  X"40",
  X"40",  X"00",  X"80",  X"00",  X"A0",  X"00",  X"E2",  X"80",
  X"40",  X"60",  X"60",  X"A0",  X"60",  X"A0",  X"A0",  X"A0",
  X"A0",  X"00",  X"A0",  X"A0",  X"A0",  X"A0",  X"A0",  X"A0",
  X"A0",  X"A0",  X"00",  X"00",  X"A0",  X"60",  X"A0",  X"A0",
  X"A0",  X"A0",  X"20",  X"00",  X"00",  X"00",  X"40",  X"80",
  X"00",  X"38",  X"20",  X"E0",  X"40",  X"40",  X"A0",  X"00",
  X"00",  X"E0",  X"A0",  X"2F",  X"00",  X"00",  X"00",  X"E0",
  X"E0",  X"FF",  X"E0",  X"20",  X"E0",  X"00",  X"00",  X"20",
  X"20",  X"40",  X"40",  X"E0",  X"00",  X"00",  X"20",  X"E0",
  X"2F",  X"00",  X"00",  X"00",  X"20",  X"20",  X"FF",  X"20",
  X"20",  X"E0",  X"00",  X"20",  X"FC",  X"40",  X"80",  X"20",
  X"40",  X"00",  X"23",  X"80",  X"A0",  X"80",  X"40",  X"E0",
  X"00",  X"00",  X"E0",  X"62",  X"BF",  X"00",  X"20",  X"3F",
  X"7F",  X"00",  X"3F",  X"40",  X"3F",  X"00",  X"7F",  X"FF",
  X"00",  X"E0",  X"00",  X"BF",  X"E0",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"52",  X"0F",  X"0E",  X"00",  X"00",  X"6D",
  X"00",  X"00",  X"00",  X"00",  X"50",  X"7C",  X"40",  X"1B",
  X"00",  X"00",  X"00",  X"6C",  X"00",  X"0D",  X"09",  X"00",
  X"00",  X"00",  X"6D",  X"00",  X"0D",  X"09",  X"00",  X"00",
  X"00",  X"6D",  X"01",  X"0D",  X"09",  X"00",  X"00",  X"00",
  X"6E",  X"01",  X"0D",  X"09",  X"00",  X"00",  X"00",  X"6F",
  X"00",  X"0D",  X"09",  X"00",  X"00",  X"00",  X"6F",  X"00",
  X"0D",  X"09",  X"00",  X"00",  X"00",  X"70",  X"00",  X"0D",
  X"09",  X"00",  X"00",  X"00",  X"70",  X"00",  X"0D",  X"09",
  X"00",  X"00",  X"01",  X"71",  X"00",  X"0D",  X"09",  X"00",
  X"00",  X"01",  X"71",  X"00",  X"0D",  X"09",  X"00",  X"00",
  X"01",  X"71",  X"00",  X"0D",  X"09",  X"00",  X"00",  X"01",
  X"71",  X"00",  X"00",  X"00",  X"01",  X"71",  X"00",  X"0D",
  X"09",  X"00",  X"00",  X"01",  X"71",  X"00",  X"0D",  X"09",
  X"00",  X"00",  X"01",  X"72",  X"01",  X"0D",  X"09",  X"00",
  X"00",  X"01",  X"73",  X"00",  X"00",  X"00",  X"01",  X"73",
  X"00",  X"00",  X"00",  X"02",  X"73",  X"06",  X"0D",  X"09",
  X"00",  X"00",  X"02",  X"7A",  X"00",  X"00",  X"00",  X"02",
  X"7A",  X"00",  X"00",  X"00",  X"02",  X"7A",  X"00",  X"0D",
  X"09",  X"00",  X"00",  X"02",  X"7B",  X"00",  X"0D",  X"09",
  X"00",  X"00",  X"02",  X"7B",  X"1D",  X"0D",  X"0F",  X"00",
  X"02",  X"98",  X"00",  X"00",  X"00",  X"02",  X"99",  X"00",
  X"0D",  X"09",  X"00",  X"00",  X"02",  X"99",  X"00",  X"00",
  X"00",  X"02",  X"99",  X"01",  X"0D",  X"09",  X"00",  X"00",
  X"03",  X"9A",  X"00",  X"00",  X"00",  X"03",  X"9A",  X"03",
  X"0D",  X"09",  X"00",  X"00",  X"03",  X"9E",  X"01",  X"0D",
  X"09",  X"00",  X"00",  X"03",  X"9F",  X"02",  X"0D",  X"09",
  X"00",  X"00",  X"03",  X"A1",  X"13",  X"0D",  X"09",  X"00",
  X"00",  X"03",  X"B4",  X"01",  X"0D",  X"09",  X"00",  X"00",
  X"03",  X"B5",  X"00",  X"00",  X"00",  X"03",  X"B5",  X"00",
  X"00",  X"00",  X"03",  X"B5",  X"00",  X"0D",  X"09",  X"00",
  X"00",  X"03",  X"B5",  X"00",  X"00",  X"00",  X"03",  X"B5",
  X"00",  X"0D",  X"09",  X"00",  X"00",  X"04",  X"B5",  X"00",
  X"0D",  X"09",  X"00",  X"00",  X"04",  X"B5",  X"00",  X"00",
  X"00",  X"04",  X"B5",  X"00",  X"0D",  X"0F",  X"00",  X"04",
  X"B5",  X"00",  X"0D",  X"09",  X"00",  X"00",  X"04",  X"B6",
  X"00",  X"0D",  X"09",  X"00",  X"00",  X"04",  X"B6",  X"00",
  X"0D",  X"09",  X"00",  X"00",  X"04",  X"B6",  X"01",  X"0D",
  X"0F",  X"00",  X"04",  X"B7",  X"00",  X"0D",  X"0F",  X"00",
  X"04",  X"B8",  X"02",  X"0D",  X"09",  X"00",  X"00",  X"04",
  X"BB",  X"04",  X"0D",  X"09",  X"00",  X"00",  X"05",  X"BF",
  X"00",  X"0D",  X"0F",  X"00",  X"05",  X"BF",  X"00",  X"0D",
  X"0F",  X"00",  X"05",  X"C0",  X"00",  X"00",  X"00",  X"05",
  X"C0",  X"00",  X"00",  X"00",  X"05",  X"C0",  X"00",  X"00",
  X"00",  X"05",  X"C0",  X"00",  X"0D",  X"09",  X"00",  X"00",
  X"05",  X"C0",  X"00",  X"00",  X"00",  X"05",  X"C1",  X"01",
  X"0D",  X"09",  X"00",  X"00",  X"05",  X"C2",  X"00",  X"0D",
  X"09",  X"00",  X"00",  X"05",  X"C3",  X"00",  X"0D",  X"09",
  X"00",  X"00",  X"06",  X"C4",  X"01",  X"0D",  X"09",  X"00",
  X"00",  X"06",  X"C5",  X"00",  X"0D",  X"09",  X"00",  X"00",
  X"06",  X"C5",  X"00",  X"00",  X"00",  X"06",  X"C6",  X"00",
  X"00",  X"00",  X"06",  X"C6",  X"00",  X"00",  X"00",  X"06",
  X"C7",  X"00",  X"0D",  X"09",  X"00",  X"00",  X"06",  X"C7",
  X"00",  X"0E",  X"00",  X"06",  X"C8",  X"01",  X"0D",  X"09",
  X"00",  X"00",  X"06",  X"C9",  X"00",  X"0D",  X"09",  X"00",
  X"00",  X"06",  X"C9",  X"00",  X"00",  X"00",  X"06",  X"C9",
  X"00",  X"0D",  X"09",  X"00",  X"00",  X"07",  X"CA",  X"01",
  X"0D",  X"09",  X"00",  X"00",  X"07",  X"CB",  X"01",  X"0D",
  X"09",  X"00",  X"00",  X"07",  X"CD",  X"01",  X"0D",  X"09",
  X"00",  X"00",  X"07",  X"CE",  X"02",  X"0D",  X"09",  X"00",
  X"00",  X"07",  X"D0",  X"00",  X"0D",  X"09",  X"00",  X"00",
  X"07",  X"D0",  X"00",  X"0D",  X"09",  X"00",  X"00",  X"07",
  X"D1",  X"01",  X"0D",  X"09",  X"00",  X"00",  X"07",  X"D1",
  X"00",  X"0D",  X"09",  X"00",  X"00",  X"07",  X"D2",  X"04",
  X"0D",  X"09",  X"00",  X"00",  X"08",  X"D7",  X"00",  X"0D",
  X"09",  X"00",  X"00",  X"08",  X"D7",  X"00",  X"0D",  X"09",
  X"00",  X"00",  X"08",  X"D8",  X"01",  X"0D",  X"09",  X"00",
  X"00",  X"08",  X"D8",  X"00",  X"00",  X"00",  X"08",  X"D9",
  X"00",  X"00",  X"00",  X"08",  X"D9",  X"00",  X"00",  X"00",
  X"08",  X"D9",  X"00",  X"0D",  X"09",  X"00",  X"00",  X"08",
  X"D9",  X"00",  X"0D",  X"09",  X"00",  X"00",  X"08",  X"D9",
  X"00",  X"0D",  X"09",  X"00",  X"00",  X"08",  X"D9",  X"00",
  X"00",  X"00",  X"09",  X"DA",  X"00",  X"0D",  X"09",  X"00",
  X"00",  X"09",  X"DB",  X"00",  X"0D",  X"09",  X"00",  X"00",
  X"09",  X"DB",  X"00",  X"0D",  X"09",  X"00",  X"00",  X"09",
  X"DB",  X"00",  X"0D",  X"09",  X"00",  X"00",  X"09",  X"DB",
  X"01",  X"0D",  X"09",  X"00",  X"00",  X"09",  X"DD",  X"00",
  X"00",  X"00",  X"09",  X"DD",  X"00",  X"0D",  X"09",  X"00",
  X"00",  X"09",  X"DD",  X"00",  X"0D",  X"09",  X"00",  X"00",
  X"09",  X"DD",  X"00",  X"0D",  X"09",  X"00",  X"00",  X"09",
  X"E4",  X"00",  X"00",  X"00",  X"0A",  X"E4",  X"00",  X"00",
  X"00",  X"0A",  X"E4",  X"00",  X"00",  X"00",  X"0A",  X"E4",
  X"00",  X"0D",  X"0F",  X"00",  X"0A",  X"E4",  X"00",  X"0D",
  X"09",  X"00",  X"00",  X"0A",  X"E4",  X"00",  X"00",  X"00",
  X"0A",  X"E4",  X"00",  X"0D",  X"09",  X"00",  X"00",  X"0A",
  X"E4",  X"00",  X"00",  X"00",  X"0A",  X"E5",  X"00",  X"00",
  X"00",  X"0A",  X"E9",  X"00",  X"0D",  X"09",  X"00",  X"00",
  X"0A",  X"EA",  X"00",  X"00",  X"00",  X"0A",  X"EA",  X"01",
  X"0D",  X"09",  X"00",  X"00",  X"0B",  X"EC",  X"00",  X"00",
  X"00",  X"0B",  X"EC",  X"00",  X"0D",  X"09",  X"00",  X"00",
  X"0B",  X"EC",  X"00",  X"0D",  X"09",  X"00",  X"00",  X"0B",
  X"EC",  X"00",  X"0D",  X"09",  X"00",  X"00",  X"0B",  X"EC",
  X"00",  X"0D",  X"09",  X"00",  X"00",  X"0B",  X"EC",  X"00",
  X"0D",  X"09",  X"00",  X"00",  X"0B",  X"EC",  X"00",  X"0D",
  X"09",  X"00",  X"00",  X"0B",  X"ED",  X"00",  X"0D",  X"09",
  X"00",  X"00",  X"0B",  X"ED",  X"00",  X"0D",  X"09",  X"00",
  X"00",  X"0C",  X"EE",  X"00",  X"0D",  X"09",  X"00",  X"00",
  X"0C",  X"F3",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"FF",  X"00",  X"00",  X"00",  X"FF",  X"00",  X"00",
  X"01",  X"02",  X"03",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"01",  X"02",  X"04",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"01",  X"02",
  X"04",  X"08",  X"10",  X"20",  X"40",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"01",  X"02",  X"03",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"3A",  X"0A",  X"51",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"01",  X"02",  X"04",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"01",  X"02",  X"04",  X"08",
  X"10",  X"20",  X"40",  X"00",  X"01",  X"02",  X"03",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"01",  X"02",
  X"04",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"01",  X"02",  X"04",  X"08",  X"10",  X"20",
  X"40",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"01",  X"02",  X"04",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"01",  X"02",  X"04",
  X"08",  X"10",  X"20",  X"40",  X"01",  X"02",  X"03",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"1E",  X"85",  X"01",  X"02",
  X"03",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"01",  X"02",
  X"04",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"01",  X"02",  X"04",  X"08",  X"10",  X"20",
  X"40",  X"00",  X"B6",  X"00",  X"00",  X"00",  X"32",  X"36",
  X"41",  X"45",  X"00",  X"00",  X"66",  X"00",  X"32",  X"36",
  X"61",  X"65",  X"00",  X"00",  X"4E",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"75",  X"00",  X"00",  X"00",  X"30",  X"30",
  X"30",  X"30",  X"20",  X"20",  X"20",  X"20",  X"55",  X"38",
  X"53",  X"00",  X"45",  X"50",  X"4A",  X"00",  X"66",  X"74",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"87",  X"43",
  X"8A",  X"C8",  X"44",  X"79",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"4F",  X"35",
  X"00",  X"00",  X"B4",  X"B4",  X"B4",  X"B4",  X"B4",  X"B4",
  X"B4",  X"B4",  X"B4",  X"B4",  X"7F",  X"7F",  X"B5",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"40",  X"00",
  X"88",  X"00",  X"6A",  X"00",  X"84",  X"00",  X"12",  X"00",
  X"D7",  X"00",  X"CD",  X"00",  X"A0",  X"00",  X"48",  X"00",
  X"1A",  X"00",  X"30",  X"00",  X"BC",  X"00",  X"6B",  X"00",
  X"C3",  X"80",  X"34",  X"A0",  X"C1",  X"C8",  X"58",  X"3D",
  X"AF",  X"8C",  X"1A",  X"EF",  X"F0",  X"D5",  X"2D",  X"4A",
  X"78",  X"9D",  X"C3",  X"80",  X"B8",  X"6E",  X"4F",  X"F9",
  X"77",  X"1D",  X"4F",  X"BF",  X"D2",  X"89",  X"F6",  X"A7",
  X"0F",  X"A7",  X"BA",  X"97",  X"06",  X"6F",  X"00",  X"00",
  X"00",  X"00",  X"BF",  X"D6",  X"00",  X"FB",  X"00",  X"E0",
  X"00",  X"BF",  X"D6",  X"00",  X"E0",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"B6",  X"00",  X"00",  X"B9",
  X"BA",  X"BB",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"B4",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"AB",  X"E6",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"BC",  X"BC",  X"BC",  X"BC",
  X"BC",  X"BC",  X"BC",  X"BC",  X"BC",  X"BC",  X"BC",  X"BC",
  X"BC",  X"BC",  X"BC",  X"BC",  X"BC",  X"BC",  X"BC",  X"BC",
  X"BC",  X"BC",  X"BC",  X"BC",  X"BC",  X"BC",  X"BC",  X"BC",
  X"BC",  X"BC",  X"BC",  X"BC",  X"BC",  X"BC",  X"BC",  X"BC",
  X"BC",  X"BC",  X"BC",  X"BC",  X"BC",  X"BC",  X"BC",  X"BC",
  X"BC",  X"BC",  X"BD",  X"BD",  X"BD",  X"BD",  X"BD",  X"BD",
  X"BD",  X"BD",  X"BD",  X"BD",  X"BD",  X"BD",  X"BD",  X"BD",
  X"BD",  X"BD",  X"BD",  X"BD",  X"BD",  X"BD",  X"BD",  X"BD",
  X"BD",  X"BD",  X"BD",  X"BD",  X"BD",  X"BD",  X"BD",  X"BD",
  X"BD",  X"BD",  X"BD",  X"BD",  X"BD",  X"BD",  X"BD",  X"BD",
  X"BD",  X"BD",  X"BD",  X"BD",  X"BD",  X"BD",  X"BD",  X"BD",
  X"BD",  X"BD",  X"BD",  X"BD",  X"BD",  X"BD",  X"BD",  X"BD",
  X"BD",  X"BD",  X"BD",  X"BD",  X"BD",  X"BD",  X"BD",  X"BD",
  X"BD",  X"BD",  X"BE",  X"BE",  X"BE",  X"BE",  X"BE",  X"BE",
  X"BE",  X"BE",  X"BE",  X"BE",  X"BE",  X"BE",  X"BE",  X"BE",
  X"BE",  X"BE",  X"BE",  X"BE",  X"BE",  X"BE",  X"BE",  X"BE",
  X"BE",  X"BE",  X"BE",  X"BE",  X"BE",  X"BE",  X"BE",  X"BE",
  X"BE",  X"BE",  X"BE",  X"BE",  X"BE",  X"BE",  X"BE",  X"BE",
  X"BE",  X"BE",  X"BE",  X"BE",  X"BE",  X"BE",  X"BE",  X"BE",
  X"BE",  X"BE",  X"BE",  X"BE",  X"BE",  X"BE",  X"BE",  X"BE",
  X"BE",  X"BE",  X"BE",  X"BE",  X"BE",  X"BE",  X"BE",  X"BE",
  X"BE",  X"BE",  X"BF",  X"BF",  X"BF",  X"BF",  X"BF",  X"BF",
  X"BF",  X"BF",  X"BF",  X"BF",  X"BF",  X"BF",  X"BF",  X"BF",
  X"BF",  X"BF",  X"BF",  X"BF",  X"BF",  X"BF",  X"BF",  X"BF",
  X"BF",  X"BF",  X"BF",  X"BF",  X"BF",  X"BF",  X"BF",  X"BF",
  X"BF",  X"BF",  X"BF",  X"BF",  X"BF",  X"BF",  X"BF",  X"BF",
  X"BF",  X"BF",  X"BF",  X"BF",  X"BF",  X"BF",  X"BF",  X"BF",
  X"BF",  X"BF",  X"BF",  X"BF",  X"BF",  X"BF",  X"BF",  X"BF",
  X"BF",  X"BF",  X"BF",  X"BF",  X"BF",  X"BF",  X"BF",  X"BF",
  X"BF",  X"BF",  X"C0",  X"C0",  X"C0",  X"C0",  X"C0",  X"C0",
  X"C0",  X"C0",  X"C0",  X"C0",  X"C0",  X"C0",  X"C0",  X"C0",
  X"C0",  X"C0",  X"C0",  X"C0",  X"00",  X"FF",  X"00",  X"C0",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"C0",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"C1",  X"C1",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"01",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"8A",  X"03",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  others => X"00" );


constant ram02 : ram_type := (
  X"10",  X"10",  X"C1",  X"00",  X"48",  X"50",  X"80",  X"10",
  X"D0",  X"00",  X"00",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"48",  X"10",  X"C5",  X"00",  X"48",  X"10",  X"C5",  X"00",
  X"48",  X"10",  X"C5",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"D0",  X"00",  X"00",  X"00",  X"48",  X"50",  X"80",  X"10",
  X"D0",  X"00",  X"00",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"D0",  X"00",  X"00",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"D0",  X"00",  X"00",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"D0",  X"00",  X"00",  X"00",  X"10",  X"48",  X"80",  X"50",
  X"10",  X"48",  X"80",  X"50",  X"10",  X"48",  X"80",  X"50",
  X"10",  X"48",  X"80",  X"50",  X"10",  X"48",  X"80",  X"50",
  X"10",  X"48",  X"80",  X"50",  X"10",  X"48",  X"80",  X"50",
  X"10",  X"48",  X"80",  X"50",  X"10",  X"48",  X"80",  X"50",
  X"10",  X"48",  X"80",  X"50",  X"10",  X"48",  X"80",  X"50",
  X"10",  X"48",  X"80",  X"50",  X"10",  X"48",  X"80",  X"50",
  X"10",  X"48",  X"80",  X"50",  X"10",  X"48",  X"80",  X"50",
  X"D0",  X"00",  X"00",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"D0",  X"00",  X"00",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"D0",  X"00",  X"00",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"D0",  X"00",  X"00",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"D0",  X"00",  X"00",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"D0",  X"00",  X"00",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"D0",  X"00",  X"00",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"D0",  X"00",  X"00",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"D0",  X"00",  X"00",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"D0",  X"00",  X"00",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"D0",  X"00",  X"00",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"D0",  X"00",  X"00",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"D0",  X"00",  X"00",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"D0",  X"00",  X"00",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"D0",  X"00",  X"00",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"D0",  X"00",  X"00",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"D0",  X"00",  X"00",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"D0",  X"00",  X"00",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"D0",  X"00",  X"00",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"D0",  X"00",  X"00",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"D0",  X"00",  X"00",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"D0",  X"00",  X"00",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"D0",  X"00",  X"00",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"D0",  X"00",  X"00",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"D0",  X"00",  X"00",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"D0",  X"00",  X"00",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"D0",  X"00",  X"00",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"D0",  X"00",  X"00",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"D0",  X"00",  X"00",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"D0",  X"00",  X"00",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"D0",  X"00",  X"00",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"D0",  X"00",  X"00",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"D0",  X"00",  X"00",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"D0",  X"00",  X"00",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"D0",  X"00",  X"00",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"D0",  X"00",  X"00",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"D0",  X"00",  X"00",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"D0",  X"00",  X"00",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"D0",  X"00",  X"00",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"D0",  X"00",  X"00",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"D0",  X"00",  X"00",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"D0",  X"00",  X"00",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"D0",  X"00",  X"00",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"D0",  X"00",  X"00",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"D0",  X"00",  X"00",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"D0",  X"00",  X"00",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"D0",  X"00",  X"00",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"D0",  X"00",  X"00",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"D0",  X"00",  X"00",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"48",  X"10",  X"C5",  X"00",  X"48",  X"80",  X"50",  X"00",
  X"D0",  X"00",  X"00",  X"00",  X"48",  X"10",  X"C5",  X"00",
  X"D0",  X"00",  X"00",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"D0",  X"00",  X"00",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"D0",  X"00",  X"00",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"D0",  X"00",  X"00",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"D0",  X"00",  X"00",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"D0",  X"00",  X"00",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"D0",  X"00",  X"00",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"D0",  X"00",  X"00",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"D0",  X"00",  X"00",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"D0",  X"00",  X"00",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"D0",  X"00",  X"00",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"D0",  X"00",  X"00",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"D0",  X"00",  X"00",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"D0",  X"00",  X"00",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"D0",  X"00",  X"00",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"D0",  X"00",  X"00",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"D0",  X"00",  X"00",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"D0",  X"00",  X"00",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"D0",  X"00",  X"00",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"D0",  X"00",  X"00",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"D0",  X"00",  X"00",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"D0",  X"00",  X"00",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"D0",  X"00",  X"00",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"D0",  X"00",  X"00",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"D0",  X"00",  X"00",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"D0",  X"00",  X"00",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"D0",  X"00",  X"00",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"D0",  X"00",  X"00",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"D0",  X"00",  X"00",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"D0",  X"00",  X"00",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"D0",  X"00",  X"00",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"D0",  X"00",  X"00",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"D0",  X"00",  X"00",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"D0",  X"00",  X"00",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"D0",  X"00",  X"00",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"D0",  X"00",  X"00",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"D0",  X"00",  X"00",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"D0",  X"00",  X"00",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"D0",  X"00",  X"00",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"D0",  X"00",  X"00",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"D0",  X"00",  X"00",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"D0",  X"00",  X"00",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"D0",  X"00",  X"00",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"D0",  X"00",  X"00",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"D0",  X"00",  X"00",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"D0",  X"00",  X"00",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"D0",  X"00",  X"00",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"D0",  X"00",  X"00",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"D0",  X"00",  X"00",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"D0",  X"00",  X"00",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"D0",  X"00",  X"00",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"D0",  X"00",  X"00",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"D0",  X"00",  X"00",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"D0",  X"00",  X"00",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"D0",  X"00",  X"00",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"D0",  X"00",  X"00",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"D0",  X"00",  X"00",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"D0",  X"00",  X"00",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"D0",  X"00",  X"00",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"D0",  X"00",  X"00",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"D0",  X"00",  X"00",  X"00",  X"D0",  X"00",  X"00",  X"00",
  X"E3",  X"10",  X"10",  X"10",  X"10",  X"10",  X"20",  X"A0",
  X"BF",  X"38",  X"10",  X"12",  X"22",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"10",  X"12",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"C7",  X"E8",  X"E3",
  X"10",  X"0C",  X"A0",  X"80",  X"10",  X"04",  X"10",  X"10",
  X"14",  X"14",  X"24",  X"3C",  X"04",  X"A0",  X"80",  X"00",
  X"14",  X"00",  X"28",  X"24",  X"04",  X"C0",  X"00",  X"04",
  X"A0",  X"BF",  X"00",  X"00",  X"10",  X"A0",  X"80",  X"10",
  X"10",  X"FF",  X"12",  X"10",  X"2C",  X"C7",  X"E8",  X"E3",
  X"C7",  X"E8",  X"E3",  X"00",  X"10",  X"A0",  X"80",  X"10",
  X"10",  X"10",  X"12",  X"FF",  X"12",  X"10",  X"02",  X"A0",
  X"80",  X"12",  X"00",  X"10",  X"A0",  X"80",  X"00",  X"C0",
  X"00",  X"C7",  X"E8",  X"E3",  X"C7",  X"E8",  X"C3",  X"00",
  X"E3",  X"27",  X"27",  X"27",  X"27",  X"27",  X"27",  X"27",
  X"07",  X"27",  X"07",  X"10",  X"10",  X"07",  X"10",  X"00",
  X"00",  X"10",  X"27",  X"10",  X"10",  X"10",  X"10",  X"07",
  X"00",  X"00",  X"07",  X"10",  X"E8",  X"C3",  X"00",  X"E3",
  X"10",  X"10",  X"00",  X"00",  X"E8",  X"C3",  X"00",  X"E3",
  X"27",  X"07",  X"00",  X"A0",  X"80",  X"00",  X"07",  X"00",
  X"07",  X"00",  X"00",  X"3F",  X"10",  X"08",  X"20",  X"80",
  X"00",  X"07",  X"00",  X"07",  X"00",  X"07",  X"00",  X"20",
  X"00",  X"08",  X"28",  X"38",  X"20",  X"07",  X"00",  X"00",
  X"07",  X"20",  X"07",  X"00",  X"18",  X"A0",  X"60",  X"08",
  X"A0",  X"80",  X"00",  X"07",  X"00",  X"07",  X"00",  X"00",
  X"3F",  X"10",  X"08",  X"20",  X"80",  X"00",  X"07",  X"00",
  X"00",  X"08",  X"18",  X"A0",  X"60",  X"08",  X"A0",  X"BF",
  X"00",  X"E8",  X"C3",  X"00",  X"E3",  X"27",  X"27",  X"27",
  X"07",  X"27",  X"07",  X"00",  X"07",  X"00",  X"07",  X"20",
  X"07",  X"00",  X"A0",  X"80",  X"00",  X"07",  X"10",  X"20",
  X"27",  X"80",  X"00",  X"07",  X"00",  X"07",  X"00",  X"00",
  X"07",  X"07",  X"01",  X"08",  X"28",  X"08",  X"28",  X"07",
  X"00",  X"00",  X"07",  X"20",  X"07",  X"00",  X"07",  X"00",
  X"A0",  X"60",  X"08",  X"A0",  X"80",  X"00",  X"07",  X"00",
  X"07",  X"20",  X"07",  X"00",  X"27",  X"10",  X"07",  X"07",
  X"A0",  X"80",  X"00",  X"10",  X"08",  X"A0",  X"BF",  X"00",
  X"07",  X"00",  X"A0",  X"80",  X"00",  X"07",  X"00",  X"07",
  X"00",  X"00",  X"10",  X"00",  X"10",  X"20",  X"07",  X"FF",
  X"00",  X"E8",  X"C3",  X"00",  X"E3",  X"27",  X"07",  X"20",
  X"10",  X"20",  X"07",  X"00",  X"10",  X"20",  X"07",  X"00",
  X"07",  X"20",  X"07",  X"20",  X"07",  X"00",  X"00",  X"10",
  X"20",  X"E8",  X"C3",  X"00",  X"E3",  X"27",  X"07",  X"20",
  X"10",  X"20",  X"07",  X"00",  X"10",  X"20",  X"07",  X"00",
  X"10",  X"20",  X"27",  X"80",  X"00",  X"07",  X"00",  X"07",
  X"28",  X"00",  X"20",  X"07",  X"00",  X"27",  X"10",  X"07",
  X"A0",  X"80",  X"00",  X"10",  X"08",  X"A0",  X"BF",  X"00",
  X"07",  X"00",  X"00",  X"10",  X"20",  X"07",  X"00",  X"10",
  X"20",  X"E8",  X"C3",  X"00",  X"E3",  X"10",  X"10",  X"00",
  X"00",  X"10",  X"10",  X"20",  X"10",  X"10",  X"00",  X"10",
  X"10",  X"10",  X"10",  X"10",  X"FF",  X"00",  X"E8",  X"C3",
  X"00",  X"E3",  X"27",  X"07",  X"20",  X"10",  X"20",  X"07",
  X"00",  X"20",  X"07",  X"00",  X"20",  X"07",  X"00",  X"10",
  X"20",  X"10",  X"10",  X"10",  X"00",  X"00",  X"10",  X"10",
  X"10",  X"00",  X"00",  X"07",  X"00",  X"07",  X"00",  X"00",
  X"10",  X"20",  X"07",  X"00",  X"07",  X"00",  X"00",  X"10",
  X"20",  X"E8",  X"C3",  X"00",  X"E3",  X"27",  X"27",  X"07",
  X"00",  X"07",  X"00",  X"00",  X"10",  X"07",  X"29",  X"38",
  X"08",  X"20",  X"E8",  X"C3",  X"00",  X"E3",  X"27",  X"10",
  X"10",  X"FF",  X"00",  X"07",  X"00",  X"10",  X"FF",  X"00",
  X"07",  X"10",  X"FF",  X"00",  X"E8",  X"C3",  X"00",  X"E3",
  X"10",  X"10",  X"FF",  X"00",  X"10",  X"10",  X"18",  X"3F",
  X"10",  X"27",  X"80",  X"00",  X"10",  X"10",  X"10",  X"10",
  X"13",  X"00",  X"10",  X"00",  X"E3",  X"10",  X"37",  X"1F",
  X"10",  X"27",  X"27",  X"10",  X"27",  X"37",  X"10",  X"27",
  X"10",  X"10",  X"00",  X"07",  X"07",  X"28",  X"C7",  X"E8",
  X"E3",  X"10",  X"00",  X"10",  X"37",  X"1F",  X"10",  X"27",
  X"27",  X"10",  X"27",  X"27",  X"37",  X"10",  X"10",  X"00",
  X"07",  X"07",  X"28",  X"C7",  X"E8",  X"E3",  X"10",  X"00",
  X"14",  X"10",  X"00",  X"04",  X"A2",  X"80",  X"04",  X"02",
  X"A0",  X"80",  X"00",  X"A6",  X"80",  X"00",  X"02",  X"00",
  X"00",  X"28",  X"28",  X"02",  X"22",  X"22",  X"10",  X"28",
  X"10",  X"22",  X"A6",  X"80",  X"10",  X"00",  X"28",  X"00",
  X"22",  X"22",  X"10",  X"00",  X"14",  X"C7",  X"E8",  X"00",
  X"10",  X"A2",  X"80",  X"14",  X"04",  X"22",  X"24",  X"22",
  X"22",  X"22",  X"BF",  X"10",  X"02",  X"10",  X"10",  X"00",
  X"28",  X"22",  X"00",  X"22",  X"22",  X"10",  X"00",  X"14",
  X"C7",  X"E8",  X"BF",  X"24",  X"00",  X"10",  X"C7",  X"E8",
  X"10",  X"10",  X"00",  X"13",  X"00",  X"10",  X"00",  X"10",
  X"10",  X"00",  X"13",  X"00",  X"10",  X"00",  X"E3",  X"10",
  X"06",  X"A0",  X"80",  X"10",  X"08",  X"34",  X"A4",  X"80",
  X"88",  X"80",  X"00",  X"00",  X"10",  X"A4",  X"80",  X"34",
  X"10",  X"14",  X"04",  X"00",  X"A4",  X"80",  X"34",  X"04",
  X"04",  X"04",  X"08",  X"04",  X"00",  X"11",  X"20",  X"20",
  X"20",  X"10",  X"00",  X"04",  X"C7",  X"E8",  X"04",  X"04",
  X"0D",  X"25",  X"A0",  X"80",  X"A4",  X"10",  X"10",  X"00",
  X"05",  X"05",  X"A0",  X"80",  X"05",  X"05",  X"0D",  X"10",
  X"00",  X"10",  X"A2",  X"80",  X"10",  X"04",  X"A0",  X"80",
  X"10",  X"A4",  X"80",  X"05",  X"04",  X"00",  X"08",  X"20",
  X"A0",  X"80",  X"A4",  X"00",  X"10",  X"C7",  X"E8",  X"34",
  X"A0",  X"80",  X"2B",  X"A0",  X"80",  X"34",  X"00",  X"A0",
  X"80",  X"2B",  X"A0",  X"80",  X"A0",  X"34",  X"03",  X"2B",
  X"10",  X"14",  X"04",  X"00",  X"A0",  X"80",  X"04",  X"80",
  X"03",  X"80",  X"04",  X"04",  X"A0",  X"80",  X"03",  X"04",
  X"08",  X"20",  X"A0",  X"BF",  X"A0",  X"03",  X"03",  X"10",
  X"10",  X"00",  X"A0",  X"80",  X"04",  X"04",  X"08",  X"20",
  X"A0",  X"80",  X"A0",  X"20",  X"80",  X"20",  X"A0",  X"80",
  X"30",  X"30",  X"A0",  X"80",  X"00",  X"30",  X"01",  X"29",
  X"04",  X"03",  X"A0",  X"80",  X"00",  X"80",  X"04",  X"A3",
  X"80",  X"00",  X"00",  X"09",  X"A0",  X"BF",  X"00",  X"00",
  X"24",  X"24",  X"20",  X"20",  X"04",  X"3B",  X"10",  X"29",
  X"A0",  X"BF",  X"04",  X"88",  X"80",  X"0B",  X"2B",  X"10",
  X"04",  X"10",  X"03",  X"A3",  X"80",  X"04",  X"80",  X"02",
  X"80",  X"04",  X"04",  X"A3",  X"80",  X"02",  X"04",  X"08",
  X"20",  X"A0",  X"BF",  X"A0",  X"04",  X"04",  X"04",  X"14",
  X"23",  X"21",  X"20",  X"20",  X"24",  X"20",  X"20",  X"80",
  X"20",  X"04",  X"04",  X"00",  X"11",  X"20",  X"20",  X"20",
  X"10",  X"00",  X"04",  X"C7",  X"E8",  X"04",  X"00",  X"10",
  X"20",  X"10",  X"00",  X"04",  X"C7",  X"E8",  X"03",  X"BF",
  X"2B",  X"28",  X"04",  X"01",  X"04",  X"24",  X"24",  X"38",
  X"10",  X"23",  X"28",  X"21",  X"10",  X"BF",  X"24",  X"29",
  X"88",  X"BF",  X"03",  X"BF",  X"2B",  X"BF",  X"10",  X"04",
  X"04",  X"14",  X"10",  X"24",  X"20",  X"10",  X"24",  X"00",
  X"04",  X"C7",  X"E8",  X"04",  X"BF",  X"14",  X"8A",  X"BF",
  X"04",  X"8B",  X"80",  X"02",  X"00",  X"A2",  X"BF",  X"03",
  X"04",  X"29",  X"A1",  X"BF",  X"A1",  X"BF",  X"04",  X"89",
  X"80",  X"29",  X"BF",  X"10",  X"04",  X"00",  X"A0",  X"BF",
  X"03",  X"BF",  X"04",  X"05",  X"05",  X"A0",  X"80",  X"25",
  X"05",  X"A0",  X"80",  X"10",  X"04",  X"20",  X"25",  X"8C",
  X"80",  X"00",  X"10",  X"20",  X"04",  X"20",  X"04",  X"10",
  X"0D",  X"20",  X"00",  X"10",  X"A2",  X"80",  X"10",  X"22",
  X"00",  X"10",  X"05",  X"05",  X"25",  X"24",  X"A4",  X"80",
  X"24",  X"A5",  X"80",  X"05",  X"08",  X"04",  X"04",  X"09",
  X"10",  X"24",  X"10",  X"20",  X"A0",  X"80",  X"20",  X"10",
  X"00",  X"A0",  X"80",  X"20",  X"10",  X"00",  X"A0",  X"BF",
  X"20",  X"BF",  X"04",  X"BF",  X"04",  X"BF",  X"80",  X"A0",
  X"34",  X"03",  X"BF",  X"2B",  X"A0",  X"BF",  X"29",  X"A0",
  X"80",  X"A0",  X"30",  X"01",  X"BF",  X"29",  X"39",  X"10",
  X"28",  X"13",  X"24",  X"BF",  X"10",  X"10",  X"BF",  X"10",
  X"34",  X"03",  X"BF",  X"2B",  X"10",  X"BF",  X"24",  X"80",
  X"A0",  X"30",  X"01",  X"BF",  X"29",  X"88",  X"BF",  X"05",
  X"04",  X"05",  X"10",  X"BF",  X"20",  X"BF",  X"20",  X"04",
  X"00",  X"10",  X"10",  X"BF",  X"00",  X"BF",  X"10",  X"10",
  X"BF",  X"10",  X"30",  X"01",  X"BF",  X"29",  X"04",  X"28",
  X"BF",  X"24",  X"BF",  X"02",  X"10",  X"12",  X"13",  X"00",
  X"10",  X"00",  X"10",  X"12",  X"13",  X"00",  X"10",  X"00",
  X"E3",  X"10",  X"10",  X"00",  X"24",  X"A2",  X"80",  X"04",
  X"C7",  X"E8",  X"A0",  X"BF",  X"00",  X"26",  X"C7",  X"E8",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"E3",  X"06",  X"A0",  X"80",  X"10",  X"26",  X"C7",
  X"E8",  X"00",  X"10",  X"26",  X"26",  X"C7",  X"E8",  X"E3",
  X"00",  X"00",  X"02",  X"16",  X"27",  X"88",  X"80",  X"27",
  X"10",  X"00",  X"A2",  X"80",  X"16",  X"02",  X"A0",  X"80",
  X"00",  X"16",  X"88",  X"80",  X"10",  X"06",  X"A0",  X"80",
  X"08",  X"A0",  X"80",  X"56",  X"07",  X"27",  X"27",  X"27",
  X"27",  X"27",  X"27",  X"27",  X"10",  X"10",  X"14",  X"14",
  X"10",  X"10",  X"4E",  X"A0",  X"80",  X"0E",  X"A0",  X"80",
  X"28",  X"10",  X"05",  X"4D",  X"A0",  X"80",  X"A0",  X"BF",
  X"05",  X"A5",  X"80",  X"10",  X"24",  X"24",  X"04",  X"07",
  X"07",  X"00",  X"00",  X"27",  X"A0",  X"80",  X"27",  X"0D",
  X"10",  X"06",  X"28",  X"A0",  X"80",  X"06",  X"2F",  X"10",
  X"0E",  X"2D",  X"10",  X"10",  X"10",  X"10",  X"3D",  X"06",
  X"05",  X"A0",  X"80",  X"28",  X"A5",  X"80",  X"10",  X"2F",
  X"2F",  X"27",  X"27",  X"10",  X"07",  X"10",  X"8D",  X"80",
  X"8D",  X"07",  X"00",  X"27",  X"80",  X"27",  X"4F",  X"A0",
  X"80",  X"8D",  X"10",  X"24",  X"07",  X"24",  X"07",  X"07",
  X"00",  X"00",  X"27",  X"27",  X"A0",  X"80",  X"04",  X"07",
  X"A0",  X"80",  X"07",  X"07",  X"20",  X"A0",  X"80",  X"A0",
  X"80",  X"27",  X"10",  X"10",  X"10",  X"80",  X"10",  X"04",
  X"A4",  X"80",  X"10",  X"20",  X"20",  X"00",  X"07",  X"07",
  X"00",  X"01",  X"27",  X"A0",  X"BF",  X"27",  X"27",  X"10",
  X"FF",  X"07",  X"A2",  X"80",  X"07",  X"04",  X"A4",  X"BF",
  X"10",  X"10",  X"10",  X"10",  X"24",  X"07",  X"24",  X"07",
  X"00",  X"27",  X"07",  X"00",  X"27",  X"A0",  X"80",  X"04",
  X"10",  X"FF",  X"07",  X"A2",  X"80",  X"10",  X"8D",  X"80",
  X"A5",  X"24",  X"24",  X"04",  X"07",  X"00",  X"27",  X"07",
  X"00",  X"A0",  X"80",  X"27",  X"8D",  X"80",  X"07",  X"07",
  X"27",  X"A5",  X"80",  X"A5",  X"80",  X"27",  X"10",  X"80",
  X"07",  X"05",  X"A5",  X"80",  X"24",  X"24",  X"24",  X"04",
  X"07",  X"07",  X"00",  X"00",  X"27",  X"A0",  X"BF",  X"27",
  X"10",  X"FF",  X"10",  X"A2",  X"80",  X"05",  X"A5",  X"BF",
  X"10",  X"24",  X"07",  X"24",  X"07",  X"05",  X"07",  X"00",
  X"27",  X"A0",  X"80",  X"27",  X"10",  X"FF",  X"07",  X"A2",
  X"80",  X"A5",  X"07",  X"07",  X"A7",  X"80",  X"10",  X"A5",
  X"80",  X"06",  X"27",  X"A5",  X"BF",  X"10",  X"07",  X"00",
  X"10",  X"BF",  X"4E",  X"10",  X"10",  X"00",  X"C0",  X"00",
  X"BF",  X"0D",  X"15",  X"8D",  X"80",  X"06",  X"8D",  X"80",
  X"06",  X"16",  X"A0",  X"06",  X"40",  X"10",  X"2F",  X"A5",
  X"80",  X"0D",  X"07",  X"A5",  X"80",  X"27",  X"88",  X"80",
  X"88",  X"08",  X"A0",  X"80",  X"A0",  X"80",  X"07",  X"0F",
  X"05",  X"00",  X"37",  X"A7",  X"BF",  X"2D",  X"07",  X"8D",
  X"80",  X"20",  X"A0",  X"80",  X"10",  X"05",  X"20",  X"80",
  X"2D",  X"A0",  X"06",  X"40",  X"BF",  X"10",  X"15",  X"8D",
  X"80",  X"06",  X"8D",  X"80",  X"06",  X"16",  X"A0",  X"06",
  X"40",  X"BF",  X"10",  X"A0",  X"06",  X"40",  X"BF",  X"10",
  X"15",  X"8D",  X"80",  X"8D",  X"06",  X"06",  X"A7",  X"80",
  X"A0",  X"10",  X"BF",  X"40",  X"80",  X"07",  X"8D",  X"80",
  X"10",  X"07",  X"10",  X"A7",  X"80",  X"27",  X"27",  X"27",
  X"10",  X"4F",  X"A0",  X"BF",  X"8D",  X"07",  X"00",  X"27",
  X"8D",  X"BF",  X"27",  X"07",  X"27",  X"A0",  X"BF",  X"A0",
  X"80",  X"27",  X"10",  X"10",  X"10",  X"80",  X"10",  X"04",
  X"A4",  X"80",  X"10",  X"20",  X"20",  X"00",  X"07",  X"07",
  X"00",  X"01",  X"27",  X"A0",  X"BF",  X"27",  X"27",  X"10",
  X"FF",  X"07",  X"A2",  X"80",  X"07",  X"04",  X"A4",  X"BF",
  X"10",  X"10",  X"10",  X"10",  X"24",  X"07",  X"24",  X"07",
  X"00",  X"27",  X"07",  X"00",  X"27",  X"A0",  X"BF",  X"04",
  X"10",  X"FF",  X"07",  X"A2",  X"80",  X"4F",  X"A0",  X"BF",
  X"10",  X"8D",  X"BF",  X"07",  X"2F",  X"10",  X"2F",  X"10",
  X"24",  X"07",  X"24",  X"07",  X"07",  X"00",  X"00",  X"27",
  X"27",  X"A0",  X"BF",  X"04",  X"10",  X"FF",  X"07",  X"A2",
  X"80",  X"07",  X"A0",  X"BF",  X"10",  X"07",  X"27",  X"A0",
  X"BF",  X"A0",  X"80",  X"27",  X"10",  X"10",  X"10",  X"80",
  X"10",  X"04",  X"A4",  X"80",  X"10",  X"20",  X"20",  X"00",
  X"07",  X"07",  X"00",  X"01",  X"27",  X"A0",  X"BF",  X"27",
  X"27",  X"10",  X"FF",  X"07",  X"A2",  X"80",  X"07",  X"04",
  X"A4",  X"BF",  X"10",  X"10",  X"10",  X"10",  X"24",  X"07",
  X"24",  X"07",  X"00",  X"27",  X"07",  X"00",  X"27",  X"A0",
  X"BF",  X"04",  X"10",  X"FF",  X"07",  X"A2",  X"80",  X"10",
  X"BF",  X"07",  X"80",  X"07",  X"10",  X"1F",  X"10",  X"18",
  X"AA",  X"00",  X"80",  X"07",  X"10",  X"24",  X"10",  X"10",
  X"07",  X"24",  X"07",  X"00",  X"00",  X"27",  X"27",  X"A0",
  X"80",  X"04",  X"07",  X"07",  X"A0",  X"80",  X"10",  X"8D",
  X"BF",  X"8D",  X"10",  X"24",  X"07",  X"24",  X"07",  X"07",
  X"00",  X"00",  X"27",  X"27",  X"A0",  X"80",  X"04",  X"07",
  X"00",  X"A5",  X"BF",  X"A5",  X"80",  X"27",  X"10",  X"80",
  X"07",  X"05",  X"A5",  X"80",  X"24",  X"24",  X"24",  X"04",
  X"07",  X"07",  X"00",  X"00",  X"27",  X"A0",  X"BF",  X"27",
  X"10",  X"FF",  X"10",  X"A2",  X"80",  X"10",  X"BF",  X"05",
  X"10",  X"FF",  X"07",  X"A2",  X"BF",  X"27",  X"A5",  X"80",
  X"16",  X"07",  X"00",  X"10",  X"16",  X"28",  X"30",  X"88",
  X"80",  X"00",  X"88",  X"80",  X"00",  X"C7",  X"E8",  X"C7",
  X"E8",  X"00",  X"10",  X"A2",  X"80",  X"16",  X"16",  X"10",
  X"08",  X"A0",  X"BF",  X"07",  X"56",  X"A0",  X"BF",  X"16",
  X"88",  X"80",  X"00",  X"08",  X"06",  X"27",  X"07",  X"06",
  X"27",  X"27",  X"10",  X"37",  X"37",  X"27",  X"07",  X"27",
  X"27",  X"10",  X"00",  X"27",  X"10",  X"00",  X"10",  X"10",
  X"07",  X"00",  X"10",  X"00",  X"10",  X"07",  X"07",  X"10",
  X"10",  X"FF",  X"10",  X"92",  X"80",  X"17",  X"00",  X"10",
  X"A2",  X"80",  X"10",  X"17",  X"88",  X"80",  X"00",  X"16",
  X"10",  X"36",  X"00",  X"10",  X"C7",  X"E8",  X"A0",  X"80",
  X"8D",  X"0D",  X"2F",  X"10",  X"2F",  X"10",  X"24",  X"07",
  X"24",  X"07",  X"07",  X"00",  X"00",  X"27",  X"27",  X"A0",
  X"80",  X"04",  X"10",  X"1F",  X"10",  X"18",  X"AA",  X"00",
  X"80",  X"07",  X"07",  X"00",  X"24",  X"05",  X"24",  X"07",
  X"00",  X"27",  X"07",  X"00",  X"27",  X"A0",  X"80",  X"04",
  X"07",  X"24",  X"07",  X"07",  X"24",  X"07",  X"07",  X"00",
  X"00",  X"27",  X"27",  X"A0",  X"BF",  X"04",  X"10",  X"FF",
  X"07",  X"A2",  X"BF",  X"10",  X"BF",  X"8D",  X"10",  X"FF",
  X"07",  X"A2",  X"BF",  X"10",  X"BF",  X"0D",  X"00",  X"06",
  X"BF",  X"10",  X"00",  X"00",  X"BF",  X"16",  X"00",  X"06",
  X"BF",  X"16",  X"A0",  X"80",  X"07",  X"A0",  X"80",  X"24",
  X"24",  X"07",  X"24",  X"07",  X"07",  X"00",  X"00",  X"27",
  X"27",  X"A0",  X"80",  X"04",  X"07",  X"07",  X"25",  X"A5",
  X"80",  X"A5",  X"80",  X"27",  X"10",  X"80",  X"07",  X"05",
  X"A5",  X"80",  X"24",  X"24",  X"24",  X"04",  X"07",  X"07",
  X"00",  X"00",  X"27",  X"A0",  X"BF",  X"27",  X"10",  X"FF",
  X"10",  X"A2",  X"BF",  X"10",  X"BF",  X"05",  X"07",  X"2F",
  X"BF",  X"10",  X"00",  X"A5",  X"BF",  X"A5",  X"80",  X"27",
  X"10",  X"80",  X"07",  X"05",  X"A5",  X"80",  X"24",  X"24",
  X"24",  X"04",  X"07",  X"07",  X"00",  X"00",  X"27",  X"A0",
  X"BF",  X"27",  X"10",  X"FF",  X"10",  X"A2",  X"BF",  X"10",
  X"BF",  X"05",  X"BF",  X"06",  X"56",  X"BF",  X"06",  X"00",
  X"06",  X"16",  X"BF",  X"16",  X"06",  X"A7",  X"80",  X"06",
  X"20",  X"0E",  X"15",  X"BF",  X"2D",  X"A5",  X"80",  X"8D",
  X"80",  X"07",  X"06",  X"10",  X"06",  X"07",  X"2F",  X"38",
  X"2F",  X"38",  X"27",  X"0F",  X"10",  X"BF",  X"27",  X"8D",
  X"80",  X"06",  X"8D",  X"80",  X"00",  X"06",  X"BF",  X"30",
  X"0E",  X"15",  X"BF",  X"2D",  X"0E",  X"BF",  X"2D",  X"2F",
  X"0E",  X"BF",  X"2D",  X"0E",  X"15",  X"BF",  X"2D",  X"05",
  X"10",  X"4E",  X"2F",  X"2F",  X"07",  X"00",  X"05",  X"A0",
  X"BF",  X"06",  X"BF",  X"05",  X"06",  X"A0",  X"10",  X"06",
  X"10",  X"40",  X"15",  X"27",  X"10",  X"BF",  X"10",  X"0E",
  X"15",  X"BF",  X"2D",  X"0E",  X"2D",  X"3D",  X"A0",  X"80",
  X"06",  X"BF",  X"15",  X"10",  X"10",  X"8D",  X"80",  X"27",
  X"8D",  X"80",  X"06",  X"16",  X"06",  X"A0",  X"40",  X"A0",
  X"BF",  X"10",  X"8D",  X"BF",  X"2F",  X"15",  X"BF",  X"10",
  X"4E",  X"A5",  X"80",  X"06",  X"05",  X"10",  X"A0",  X"BF",
  X"10",  X"4E",  X"28",  X"28",  X"00",  X"00",  X"05",  X"A0",
  X"BF",  X"06",  X"90",  X"BF",  X"10",  X"BF",  X"05",  X"0E",
  X"15",  X"BF",  X"2D",  X"2F",  X"06",  X"A5",  X"80",  X"06",
  X"A5",  X"80",  X"8D",  X"80",  X"27",  X"A5",  X"80",  X"10",
  X"10",  X"00",  X"10",  X"A2",  X"80",  X"27",  X"22",  X"A7",
  X"80",  X"38",  X"27",  X"10",  X"27",  X"BF",  X"10",  X"10",
  X"10",  X"8D",  X"BF",  X"27",  X"06",  X"BF",  X"06",  X"4F",
  X"A0",  X"BF",  X"0E",  X"2F",  X"0E",  X"BF",  X"2D",  X"0E",
  X"15",  X"BF",  X"2D",  X"A5",  X"80",  X"A5",  X"80",  X"A5",
  X"80",  X"A5",  X"8D",  X"80",  X"10",  X"07",  X"00",  X"10",
  X"1F",  X"3F",  X"3F",  X"06",  X"00",  X"1F",  X"A2",  X"80",
  X"10",  X"1F",  X"10",  X"18",  X"AA",  X"00",  X"80",  X"10",
  X"10",  X"10",  X"27",  X"10",  X"27",  X"15",  X"BF",  X"10",
  X"06",  X"BF",  X"20",  X"07",  X"0F",  X"08",  X"05",  X"37",
  X"A7",  X"BF",  X"2D",  X"07",  X"BF",  X"20",  X"A7",  X"80",
  X"07",  X"10",  X"10",  X"10",  X"00",  X"05",  X"02",  X"10",
  X"10",  X"00",  X"2D",  X"A2",  X"BF",  X"10",  X"10",  X"07",
  X"07",  X"00",  X"28",  X"BF",  X"20",  X"BF",  X"0D",  X"10",
  X"24",  X"24",  X"04",  X"07",  X"07",  X"00",  X"00",  X"27",
  X"A0",  X"BF",  X"27",  X"10",  X"FF",  X"07",  X"A2",  X"BF",
  X"10",  X"BF",  X"07",  X"10",  X"FF",  X"07",  X"A2",  X"BF",
  X"10",  X"BF",  X"10",  X"24",  X"07",  X"24",  X"07",  X"00",
  X"07",  X"00",  X"27",  X"27",  X"A0",  X"BF",  X"04",  X"BF",
  X"10",  X"07",  X"10",  X"10",  X"00",  X"10",  X"06",  X"07",
  X"10",  X"07",  X"00",  X"10",  X"A2",  X"80",  X"10",  X"BF",
  X"06",  X"10",  X"20",  X"2F",  X"A0",  X"10",  X"BF",  X"40",
  X"24",  X"07",  X"24",  X"07",  X"00",  X"04",  X"BF",  X"27",
  X"07",  X"00",  X"10",  X"1F",  X"3F",  X"06",  X"BF",  X"3F",
  X"27",  X"10",  X"07",  X"00",  X"10",  X"A5",  X"80",  X"10",
  X"10",  X"27",  X"10",  X"10",  X"10",  X"10",  X"80",  X"10",
  X"10",  X"07",  X"00",  X"A2",  X"80",  X"07",  X"07",  X"00",
  X"07",  X"A2",  X"80",  X"16",  X"02",  X"A0",  X"80",  X"A7",
  X"BF",  X"05",  X"10",  X"10",  X"07",  X"A7",  X"80",  X"10",
  X"27",  X"BF",  X"27",  X"24",  X"04",  X"07",  X"00",  X"27",
  X"07",  X"00",  X"A0",  X"80",  X"27",  X"10",  X"07",  X"24",
  X"10",  X"10",  X"07",  X"24",  X"07",  X"00",  X"00",  X"27",
  X"27",  X"A0",  X"80",  X"04",  X"07",  X"07",  X"20",  X"24",
  X"05",  X"24",  X"07",  X"20",  X"07",  X"BF",  X"00",  X"24",
  X"07",  X"24",  X"07",  X"00",  X"07",  X"00",  X"27",  X"27",
  X"A0",  X"80",  X"04",  X"10",  X"FF",  X"07",  X"A2",  X"BF",
  X"10",  X"8D",  X"BF",  X"8D",  X"10",  X"24",  X"10",  X"10",
  X"07",  X"24",  X"07",  X"00",  X"BF",  X"00",  X"A5",  X"BF",
  X"10",  X"BF",  X"8D",  X"10",  X"FF",  X"07",  X"A2",  X"BF",
  X"10",  X"BF",  X"07",  X"10",  X"10",  X"2F",  X"27",  X"10",
  X"15",  X"27",  X"BF",  X"10",  X"10",  X"24",  X"10",  X"10",
  X"07",  X"24",  X"07",  X"00",  X"00",  X"27",  X"27",  X"A0",
  X"80",  X"04",  X"07",  X"A0",  X"80",  X"07",  X"10",  X"24",
  X"07",  X"24",  X"07",  X"07",  X"00",  X"00",  X"27",  X"27",
  X"A0",  X"80",  X"04",  X"07",  X"20",  X"A5",  X"80",  X"A5",
  X"80",  X"27",  X"10",  X"80",  X"07",  X"05",  X"A5",  X"80",
  X"20",  X"20",  X"20",  X"00",  X"07",  X"07",  X"00",  X"00",
  X"27",  X"A0",  X"BF",  X"27",  X"10",  X"FF",  X"10",  X"A2",
  X"BF",  X"10",  X"BF",  X"05",  X"A0",  X"BF",  X"8D",  X"BF",
  X"10",  X"10",  X"FF",  X"07",  X"A2",  X"BF",  X"10",  X"BF",
  X"07",  X"10",  X"FF",  X"07",  X"A2",  X"BF",  X"10",  X"BF",
  X"07",  X"10",  X"FF",  X"07",  X"A2",  X"BF",  X"10",  X"BF",
  X"10",  X"10",  X"FF",  X"07",  X"A2",  X"BF",  X"10",  X"BF",
  X"07",  X"27",  X"00",  X"10",  X"38",  X"10",  X"38",  X"0A",
  X"BF",  X"27",  X"07",  X"A0",  X"80",  X"10",  X"27",  X"BF",
  X"16",  X"FF",  X"07",  X"A2",  X"BF",  X"16",  X"27",  X"BF",
  X"16",  X"BF",  X"10",  X"0E",  X"15",  X"BF",  X"2D",  X"00",
  X"1F",  X"A2",  X"80",  X"10",  X"15",  X"A5",  X"10",  X"80",
  X"10",  X"A5",  X"80",  X"A5",  X"80",  X"10",  X"1F",  X"3F",
  X"2F",  X"07",  X"A0",  X"80",  X"A0",  X"07",  X"07",  X"23",
  X"07",  X"07",  X"07",  X"23",  X"10",  X"00",  X"07",  X"A5",
  X"80",  X"10",  X"A5",  X"80",  X"8D",  X"10",  X"A5",  X"05",
  X"80",  X"10",  X"18",  X"1F",  X"AA",  X"00",  X"80",  X"07",
  X"27",  X"1D",  X"20",  X"A0",  X"60",  X"A5",  X"80",  X"27",
  X"A0",  X"80",  X"A5",  X"07",  X"A7",  X"80",  X"A0",  X"A5",
  X"80",  X"07",  X"A0",  X"10",  X"80",  X"10",  X"10",  X"10",
  X"07",  X"2F",  X"A7",  X"80",  X"27",  X"10",  X"2F",  X"A7",
  X"80",  X"07",  X"07",  X"10",  X"2F",  X"2F",  X"07",  X"07",
  X"A0",  X"07",  X"20",  X"07",  X"27",  X"80",  X"00",  X"07",
  X"0F",  X"88",  X"80",  X"38",  X"10",  X"27",  X"2F",  X"10",
  X"38",  X"38",  X"0F",  X"00",  X"BF",  X"27",  X"8D",  X"BF",
  X"0F",  X"BF",  X"07",  X"10",  X"FF",  X"07",  X"A2",  X"BF",
  X"10",  X"BF",  X"07",  X"27",  X"38",  X"10",  X"0F",  X"BF",
  X"27",  X"20",  X"07",  X"20",  X"07",  X"00",  X"07",  X"00",
  X"27",  X"27",  X"A0",  X"80",  X"00",  X"10",  X"FF",  X"07",
  X"A2",  X"BF",  X"10",  X"07",  X"20",  X"20",  X"00",  X"07",
  X"07",  X"00",  X"00",  X"27",  X"A0",  X"BF",  X"27",  X"BF",
  X"10",  X"10",  X"10",  X"27",  X"10",  X"15",  X"27",  X"BF",
  X"10",  X"10",  X"27",  X"10",  X"27",  X"15",  X"BF",  X"10",
  X"07",  X"FF",  X"07",  X"92",  X"80",  X"10",  X"10",  X"00",
  X"07",  X"07",  X"10",  X"07",  X"07",  X"00",  X"10",  X"A7",
  X"80",  X"38",  X"2D",  X"10",  X"38",  X"27",  X"0F",  X"BF",
  X"27",  X"88",  X"BF",  X"06",  X"00",  X"10",  X"C7",  X"E8",
  X"10",  X"10",  X"10",  X"BF",  X"07",  X"80",  X"A5",  X"80",
  X"07",  X"07",  X"A0",  X"80",  X"A7",  X"8D",  X"BF",  X"10",
  X"BF",  X"07",  X"8D",  X"BF",  X"10",  X"BF",  X"07",  X"A0",
  X"10",  X"80",  X"10",  X"28",  X"00",  X"A0",  X"BF",  X"27",
  X"BF",  X"1D",  X"07",  X"10",  X"07",  X"10",  X"00",  X"07",
  X"A2",  X"80",  X"10",  X"BF",  X"27",  X"10",  X"FF",  X"07",
  X"A2",  X"BF",  X"10",  X"BF",  X"07",  X"16",  X"10",  X"10",
  X"BF",  X"36",  X"05",  X"BF",  X"10",  X"10",  X"27",  X"10",
  X"10",  X"00",  X"05",  X"02",  X"10",  X"10",  X"00",  X"2D",
  X"07",  X"A2",  X"BF",  X"10",  X"02",  X"05",  X"10",  X"2D",
  X"A0",  X"80",  X"07",  X"BF",  X"07",  X"08",  X"00",  X"28",
  X"A0",  X"BF",  X"00",  X"BF",  X"07",  X"07",  X"BF",  X"10",
  X"A0",  X"A0",  X"10",  X"3F",  X"BF",  X"2F",  X"4D",  X"A0",
  X"80",  X"10",  X"07",  X"00",  X"BF",  X"10",  X"10",  X"80",
  X"20",  X"10",  X"07",  X"07",  X"BF",  X"10",  X"10",  X"1F",
  X"10",  X"18",  X"AA",  X"00",  X"80",  X"10",  X"10",  X"20",
  X"27",  X"BF",  X"00",  X"10",  X"20",  X"BF",  X"2F",  X"07",
  X"BF",  X"00",  X"06",  X"A5",  X"BF",  X"06",  X"0E",  X"2D",
  X"BF",  X"10",  X"A7",  X"80",  X"A5",  X"80",  X"07",  X"8D",
  X"BF",  X"0F",  X"07",  X"10",  X"BF",  X"07",  X"80",  X"05",
  X"8D",  X"BF",  X"10",  X"05",  X"BF",  X"10",  X"BF",  X"10",
  X"16",  X"10",  X"BF",  X"36",  X"10",  X"10",  X"00",  X"10",
  X"10",  X"10",  X"10",  X"13",  X"FF",  X"10",  X"00",  X"E3",
  X"A6",  X"80",  X"10",  X"10",  X"10",  X"10",  X"00",  X"10",
  X"A2",  X"80",  X"10",  X"26",  X"10",  X"24",  X"C7",  X"E8",
  X"10",  X"07",  X"10",  X"00",  X"10",  X"BF",  X"A2",  X"10",
  X"10",  X"00",  X"10",  X"10",  X"10",  X"10",  X"13",  X"FF",
  X"10",  X"00",  X"E3",  X"A6",  X"80",  X"10",  X"A6",  X"80",
  X"06",  X"04",  X"07",  X"07",  X"07",  X"10",  X"10",  X"10",
  X"FF",  X"10",  X"A2",  X"80",  X"10",  X"26",  X"A0",  X"80",
  X"27",  X"A2",  X"80",  X"27",  X"A6",  X"80",  X"06",  X"A2",
  X"80",  X"10",  X"0C",  X"2C",  X"00",  X"A2",  X"BF",  X"0C",
  X"04",  X"06",  X"00",  X"26",  X"04",  X"A0",  X"80",  X"A6",
  X"80",  X"04",  X"04",  X"07",  X"07",  X"10",  X"10",  X"FF",
  X"10",  X"A2",  X"BF",  X"26",  X"10",  X"24",  X"27",  X"C7",
  X"E8",  X"27",  X"C7",  X"E8",  X"10",  X"C7",  X"E8",  X"A6",
  X"80",  X"26",  X"27",  X"C7",  X"EE",  X"06",  X"BF",  X"10",
  X"10",  X"10",  X"10",  X"00",  X"10",  X"10",  X"10",  X"10",
  X"10",  X"13",  X"FF",  X"10",  X"00",  X"E3",  X"10",  X"00",
  X"14",  X"A2",  X"80",  X"14",  X"10",  X"00",  X"12",  X"A2",
  X"80",  X"A6",  X"80",  X"A6",  X"80",  X"2E",  X"06",  X"A0",
  X"80",  X"0E",  X"0E",  X"10",  X"3E",  X"16",  X"2E",  X"2E",
  X"C7",  X"E8",  X"14",  X"10",  X"00",  X"12",  X"A2",  X"80",
  X"A6",  X"80",  X"3E",  X"88",  X"80",  X"00",  X"2E",  X"C7",
  X"E8",  X"A6",  X"BF",  X"2E",  X"C7",  X"E8",  X"06",  X"00",
  X"10",  X"A0",  X"80",  X"3F",  X"00",  X"06",  X"10",  X"A0",
  X"80",  X"0E",  X"36",  X"11",  X"08",  X"36",  X"10",  X"08",
  X"0E",  X"10",  X"38",  X"10",  X"2E",  X"2E",  X"2E",  X"2E",
  X"C7",  X"E8",  X"3F",  X"00",  X"06",  X"10",  X"A0",  X"80",
  X"0E",  X"36",  X"13",  X"09",  X"36",  X"11",  X"08",  X"36",
  X"10",  X"08",  X"0E",  X"10",  X"38",  X"10",  X"2E",  X"2E",
  X"2E",  X"2E",  X"2E",  X"C7",  X"E8",  X"08",  X"A0",  X"80",
  X"00",  X"06",  X"08",  X"A0",  X"80",  X"10",  X"06",  X"08",
  X"A0",  X"80",  X"10",  X"2E",  X"2E",  X"C7",  X"E8",  X"14",
  X"10",  X"00",  X"12",  X"A2",  X"80",  X"A6",  X"BF",  X"3E",
  X"88",  X"BF",  X"2E",  X"00",  X"08",  X"A0",  X"80",  X"06",
  X"C7",  X"E8",  X"14",  X"10",  X"00",  X"12",  X"A2",  X"BF",
  X"A6",  X"80",  X"10",  X"3E",  X"88",  X"80",  X"10",  X"06",
  X"A0",  X"80",  X"10",  X"26",  X"2E",  X"10",  X"10",  X"2E",
  X"10",  X"2E",  X"06",  X"2E",  X"C7",  X"E8",  X"3F",  X"06",
  X"A0",  X"BF",  X"0E",  X"36",  X"10",  X"08",  X"0E",  X"10",
  X"38",  X"10",  X"2E",  X"2E",  X"2E",  X"C7",  X"E8",  X"08",
  X"A0",  X"BF",  X"06",  X"C7",  X"E8",  X"0E",  X"36",  X"13",
  X"0B",  X"36",  X"13",  X"09",  X"36",  X"11",  X"08",  X"36",
  X"10",  X"08",  X"0E",  X"10",  X"38",  X"10",  X"2E",  X"2E",
  X"2E",  X"2E",  X"2E",  X"2E",  X"C7",  X"E8",  X"00",  X"08",
  X"A0",  X"BF",  X"10",  X"06",  X"08",  X"A0",  X"80",  X"00",
  X"06",  X"A0",  X"80",  X"10",  X"10",  X"26",  X"10",  X"2E",
  X"10",  X"10",  X"2E",  X"10",  X"2E",  X"06",  X"2E",  X"2E",
  X"C7",  X"E8",  X"08",  X"A0",  X"BF",  X"10",  X"2E",  X"2E",
  X"C7",  X"E8",  X"E3",  X"10",  X"04",  X"A2",  X"80",  X"10",
  X"02",  X"A0",  X"80",  X"00",  X"14",  X"28",  X"30",  X"88",
  X"80",  X"10",  X"04",  X"A0",  X"80",  X"00",  X"14",  X"88",
  X"80",  X"88",  X"80",  X"10",  X"24",  X"10",  X"C7",  X"E8",
  X"04",  X"24",  X"C7",  X"E8",  X"04",  X"20",  X"24",  X"24",
  X"C7",  X"E8",  X"00",  X"00",  X"BF",  X"14",  X"00",  X"10",
  X"BF",  X"14",  X"88",  X"BF",  X"10",  X"88",  X"80",  X"04",
  X"10",  X"04",  X"BF",  X"34",  X"A2",  X"80",  X"08",  X"04",
  X"A2",  X"80",  X"24",  X"00",  X"04",  X"14",  X"24",  X"08",
  X"04",  X"24",  X"34",  X"10",  X"24",  X"BF",  X"34",  X"E3",
  X"06",  X"06",  X"10",  X"A4",  X"80",  X"10",  X"04",  X"2F",
  X"04",  X"06",  X"00",  X"07",  X"02",  X"10",  X"00",  X"04",
  X"07",  X"92",  X"06",  X"80",  X"04",  X"00",  X"10",  X"15",
  X"10",  X"10",  X"10",  X"05",  X"0D",  X"00",  X"10",  X"35",
  X"05",  X"00",  X"10",  X"04",  X"30",  X"08",  X"06",  X"0D",
  X"35",  X"26",  X"05",  X"38",  X"0D",  X"20",  X"00",  X"34",
  X"05",  X"34",  X"A7",  X"04",  X"35",  X"BF",  X"3E",  X"A6",
  X"80",  X"10",  X"04",  X"28",  X"04",  X"A7",  X"80",  X"24",
  X"04",  X"A0",  X"80",  X"00",  X"80",  X"24",  X"00",  X"A0",
  X"80",  X"00",  X"A7",  X"BF",  X"04",  X"24",  X"10",  X"00",
  X"10",  X"A2",  X"80",  X"00",  X"06",  X"12",  X"10",  X"10",
  X"04",  X"00",  X"33",  X"31",  X"09",  X"20",  X"0B",  X"20",
  X"00",  X"38",  X"00",  X"30",  X"04",  X"30",  X"A7",  X"00",
  X"BF",  X"38",  X"04",  X"28",  X"04",  X"00",  X"A0",  X"80",
  X"A7",  X"80",  X"24",  X"04",  X"A0",  X"80",  X"00",  X"24",
  X"C7",  X"E8",  X"00",  X"A0",  X"80",  X"24",  X"00",  X"A7",
  X"BF",  X"04",  X"24",  X"C7",  X"E8",  X"E3",  X"06",  X"27",
  X"27",  X"A0",  X"07",  X"07",  X"80",  X"1F",  X"06",  X"20",
  X"10",  X"27",  X"06",  X"28",  X"20",  X"27",  X"10",  X"00",
  X"10",  X"07",  X"26",  X"07",  X"27",  X"07",  X"A4",  X"80",
  X"10",  X"24",  X"1F",  X"0C",  X"A0",  X"80",  X"10",  X"A0",
  X"1C",  X"A0",  X"AA",  X"00",  X"80",  X"10",  X"27",  X"10",
  X"A4",  X"80",  X"16",  X"10",  X"16",  X"24",  X"C7",  X"EE",
  X"00",  X"28",  X"27",  X"10",  X"00",  X"10",  X"2C",  X"A4",
  X"10",  X"07",  X"00",  X"80",  X"27",  X"24",  X"C7",  X"E8",
  X"27",  X"00",  X"10",  X"27",  X"07",  X"A0",  X"80",  X"3F",
  X"10",  X"16",  X"A4",  X"80",  X"00",  X"4E",  X"A0",  X"80",
  X"06",  X"06",  X"24",  X"C7",  X"E8",  X"24",  X"20",  X"2C",
  X"27",  X"BF",  X"07",  X"3F",  X"27",  X"27",  X"27",  X"27",
  X"10",  X"07",  X"1F",  X"10",  X"10",  X"00",  X"07",  X"34",
  X"10",  X"89",  X"07",  X"07",  X"07",  X"80",  X"07",  X"27",
  X"07",  X"07",  X"00",  X"00",  X"20",  X"A1",  X"07",  X"80",
  X"2B",  X"00",  X"20",  X"33",  X"2C",  X"10",  X"27",  X"A0",
  X"07",  X"80",  X"A0",  X"3F",  X"01",  X"1F",  X"10",  X"3F",
  X"10",  X"03",  X"10",  X"27",  X"3F",  X"27",  X"10",  X"1B",
  X"10",  X"1F",  X"A3",  X"18",  X"A3",  X"07",  X"A0",  X"10",
  X"18",  X"A3",  X"10",  X"18",  X"A4",  X"A3",  X"1C",  X"AB",
  X"A0",  X"27",  X"00",  X"80",  X"07",  X"A0",  X"AB",  X"00",
  X"80",  X"04",  X"10",  X"A4",  X"80",  X"27",  X"2C",  X"10",
  X"10",  X"18",  X"AA",  X"00",  X"80",  X"27",  X"04",  X"00",
  X"10",  X"20",  X"A0",  X"80",  X"20",  X"10",  X"10",  X"A4",
  X"80",  X"20",  X"27",  X"27",  X"06",  X"A6",  X"80",  X"10",
  X"A6",  X"80",  X"10",  X"06",  X"10",  X"A6",  X"80",  X"10",
  X"80",  X"A6",  X"A6",  X"80",  X"A6",  X"80",  X"10",  X"10",
  X"04",  X"03",  X"91",  X"80",  X"27",  X"26",  X"A1",  X"10",
  X"80",  X"10",  X"10",  X"28",  X"00",  X"A0",  X"BF",  X"00",
  X"A5",  X"26",  X"40",  X"27",  X"08",  X"27",  X"27",  X"27",
  X"00",  X"10",  X"26",  X"10",  X"8C",  X"07",  X"07",  X"07",
  X"80",  X"07",  X"A4",  X"80",  X"07",  X"A0",  X"80",  X"10",
  X"2C",  X"A5",  X"10",  X"80",  X"18",  X"A2",  X"A5",  X"05",
  X"A0",  X"27",  X"A0",  X"A3",  X"A2",  X"07",  X"03",  X"80",
  X"2D",  X"10",  X"1B",  X"A2",  X"1C",  X"AA",  X"00",  X"80",
  X"10",  X"13",  X"80",  X"14",  X"18",  X"A2",  X"1C",  X"AA",
  X"00",  X"BF",  X"27",  X"A2",  X"00",  X"A5",  X"A0",  X"27",
  X"A0",  X"A3",  X"A2",  X"07",  X"01",  X"2C",  X"BF",  X"04",
  X"A2",  X"AB",  X"00",  X"80",  X"4C",  X"AB",  X"00",  X"BF",
  X"27",  X"27",  X"07",  X"8B",  X"80",  X"4C",  X"BF",  X"27",
  X"10",  X"AC",  X"BF",  X"16",  X"BF",  X"10",  X"3F",  X"0F",
  X"01",  X"27",  X"1F",  X"10",  X"10",  X"3F",  X"28",  X"13",
  X"BF",  X"07",  X"27",  X"10",  X"10",  X"10",  X"10",  X"10",
  X"26",  X"10",  X"27",  X"27",  X"27",  X"27",  X"00",  X"10",
  X"26",  X"10",  X"8C",  X"07",  X"07",  X"07",  X"BF",  X"07",
  X"A4",  X"80",  X"0C",  X"28",  X"10",  X"A0",  X"10",  X"A0",
  X"18",  X"3C",  X"88",  X"80",  X"10",  X"A0",  X"80",  X"A3",
  X"10",  X"10",  X"88",  X"80",  X"38",  X"18",  X"A2",  X"00",
  X"A0",  X"BF",  X"00",  X"A3",  X"07",  X"A0",  X"80",  X"27",
  X"10",  X"18",  X"AA",  X"00",  X"80",  X"00",  X"A5",  X"80",
  X"07",  X"A0",  X"80",  X"00",  X"27",  X"10",  X"1B",  X"A2",
  X"10",  X"07",  X"A0",  X"A2",  X"18",  X"A3",  X"3F",  X"3F",
  X"1F",  X"00",  X"04",  X"80",  X"27",  X"27",  X"10",  X"A5",
  X"07",  X"A0",  X"A3",  X"18",  X"A3",  X"3F",  X"3F",  X"1F",
  X"80",  X"00",  X"3F",  X"10",  X"18",  X"A2",  X"1F",  X"AA",
  X"00",  X"80",  X"27",  X"A0",  X"AA",  X"00",  X"80",  X"00",
  X"27",  X"10",  X"38",  X"07",  X"10",  X"80",  X"10",  X"A5",
  X"80",  X"A6",  X"07",  X"27",  X"27",  X"A6",  X"80",  X"07",
  X"A3",  X"80",  X"A6",  X"80",  X"10",  X"10",  X"07",  X"23",
  X"27",  X"26",  X"26",  X"07",  X"A0",  X"80",  X"A5",  X"80",
  X"A4",  X"80",  X"07",  X"27",  X"27",  X"10",  X"00",  X"10",
  X"27",  X"10",  X"10",  X"00",  X"07",  X"10",  X"10",  X"00",
  X"10",  X"07",  X"07",  X"10",  X"07",  X"A0",  X"80",  X"10",
  X"27",  X"27",  X"10",  X"00",  X"10",  X"07",  X"10",  X"A0",
  X"07",  X"80",  X"07",  X"10",  X"10",  X"00",  X"10",  X"07",
  X"07",  X"10",  X"A6",  X"80",  X"27",  X"27",  X"07",  X"A3",
  X"80",  X"10",  X"00",  X"88",  X"80",  X"10",  X"07",  X"00",
  X"27",  X"06",  X"06",  X"A6",  X"80",  X"10",  X"27",  X"27",
  X"10",  X"00",  X"10",  X"07",  X"07",  X"10",  X"A6",  X"80",
  X"10",  X"27",  X"27",  X"10",  X"00",  X"10",  X"07",  X"07",
  X"10",  X"07",  X"A1",  X"80",  X"27",  X"A5",  X"80",  X"A6",
  X"A5",  X"10",  X"80",  X"10",  X"07",  X"A3",  X"80",  X"07",
  X"27",  X"27",  X"10",  X"00",  X"10",  X"07",  X"27",  X"07",
  X"07",  X"A3",  X"80",  X"07",  X"27",  X"07",  X"10",  X"10",
  X"07",  X"08",  X"10",  X"FF",  X"10",  X"02",  X"10",  X"27",
  X"00",  X"10",  X"10",  X"27",  X"10",  X"00",  X"10",  X"02",
  X"A0",  X"10",  X"80",  X"10",  X"27",  X"10",  X"00",  X"10",
  X"07",  X"A0",  X"80",  X"07",  X"A6",  X"80",  X"A3",  X"A6",
  X"80",  X"07",  X"A3",  X"80",  X"A3",  X"80",  X"A0",  X"A6",
  X"80",  X"A0",  X"A6",  X"80",  X"A0",  X"80",  X"07",  X"A6",
  X"2C",  X"80",  X"04",  X"10",  X"10",  X"10",  X"00",  X"10",
  X"A7",  X"80",  X"10",  X"10",  X"10",  X"10",  X"00",  X"10",
  X"10",  X"10",  X"10",  X"10",  X"10",  X"00",  X"06",  X"BF",
  X"10",  X"26",  X"27",  X"BF",  X"27",  X"10",  X"18",  X"A2",
  X"08",  X"BF",  X"10",  X"80",  X"10",  X"10",  X"10",  X"27",
  X"10",  X"BF",  X"10",  X"10",  X"10",  X"10",  X"00",  X"05",
  X"10",  X"10",  X"FF",  X"10",  X"02",  X"27",  X"A5",  X"2C",
  X"10",  X"BF",  X"04",  X"07",  X"10",  X"10",  X"10",  X"00",
  X"10",  X"10",  X"00",  X"10",  X"A2",  X"80",  X"4C",  X"80",
  X"4C",  X"A0",  X"0C",  X"80",  X"04",  X"A0",  X"BF",  X"10",
  X"10",  X"2D",  X"04",  X"10",  X"00",  X"10",  X"A5",  X"BF",
  X"A7",  X"80",  X"A7",  X"80",  X"10",  X"00",  X"10",  X"10",
  X"27",  X"00",  X"10",  X"BF",  X"10",  X"80",  X"07",  X"05",
  X"A3",  X"80",  X"23",  X"07",  X"20",  X"03",  X"00",  X"27",
  X"27",  X"10",  X"26",  X"27",  X"A5",  X"80",  X"10",  X"27",
  X"10",  X"27",  X"27",  X"06",  X"06",  X"10",  X"00",  X"10",
  X"07",  X"27",  X"BF",  X"07",  X"27",  X"10",  X"A5",  X"80",
  X"A0",  X"00",  X"28",  X"10",  X"10",  X"18",  X"10",  X"18",
  X"A3",  X"A0",  X"27",  X"A0",  X"A2",  X"07",  X"00",  X"2D",
  X"3F",  X"1F",  X"A3",  X"AA",  X"00",  X"BF",  X"05",  X"10",
  X"19",  X"A3",  X"AA",  X"00",  X"80",  X"A0",  X"80",  X"10",
  X"11",  X"1B",  X"80",  X"10",  X"19",  X"A3",  X"AB",  X"00",
  X"80",  X"07",  X"80",  X"A0",  X"A3",  X"A0",  X"27",  X"A0",
  X"A3",  X"A2",  X"00",  X"AB",  X"A0",  X"07",  X"03",  X"2C",
  X"00",  X"BF",  X"04",  X"BF",  X"10",  X"07",  X"A1",  X"BF",
  X"27",  X"27",  X"3F",  X"07",  X"A8",  X"BF",  X"27",  X"1F",
  X"88",  X"BF",  X"27",  X"10",  X"06",  X"06",  X"BF",  X"27",
  X"4C",  X"A0",  X"0C",  X"BF",  X"04",  X"A0",  X"BF",  X"10",
  X"10",  X"04",  X"2D",  X"10",  X"BF",  X"10",  X"A0",  X"BF",
  X"A0",  X"10",  X"27",  X"00",  X"10",  X"07",  X"BF",  X"10",
  X"A7",  X"BF",  X"A2",  X"A5",  X"BF",  X"10",  X"18",  X"A3",
  X"AB",  X"00",  X"BF",  X"27",  X"10",  X"07",  X"10",  X"04",
  X"2D",  X"05",  X"BF",  X"10",  X"10",  X"20",  X"A0",  X"80",
  X"07",  X"00",  X"00",  X"06",  X"06",  X"BF",  X"27",  X"10",
  X"10",  X"10",  X"10",  X"00",  X"06",  X"10",  X"BF",  X"10",
  X"A0",  X"A0",  X"A0",  X"BF",  X"10",  X"08",  X"10",  X"28",
  X"10",  X"18",  X"38",  X"A2",  X"A0",  X"BF",  X"10",  X"10",
  X"10",  X"88",  X"80",  X"38",  X"18",  X"A2",  X"00",  X"A0",
  X"BF",  X"00",  X"BF",  X"07",  X"27",  X"A0",  X"A2",  X"A0",
  X"05",  X"07",  X"00",  X"10",  X"10",  X"2D",  X"3F",  X"00",
  X"28",  X"18",  X"1F",  X"80",  X"A4",  X"10",  X"1B",  X"10",
  X"A2",  X"A0",  X"27",  X"A0",  X"07",  X"01",  X"2D",  X"00",
  X"A0",  X"BF",  X"A2",  X"00",  X"04",  X"10",  X"18",  X"A4",
  X"AA",  X"00",  X"BF",  X"07",  X"A3",  X"AA",  X"00",  X"BF",
  X"00",  X"80",  X"4C",  X"10",  X"4C",  X"A0",  X"BF",  X"04",
  X"BF",  X"10",  X"10",  X"18",  X"BF",  X"A3",  X"10",  X"A7",
  X"80",  X"10",  X"27",  X"BF",  X"10",  X"BF",  X"10",  X"BF",
  X"07",  X"04",  X"00",  X"28",  X"04",  X"00",  X"27",  X"00",
  X"27",  X"10",  X"07",  X"20",  X"BF",  X"07",  X"27",  X"10",
  X"00",  X"10",  X"07",  X"A2",  X"BF",  X"07",  X"10",  X"10",
  X"10",  X"00",  X"10",  X"04",  X"10",  X"A5",  X"07",  X"07",
  X"BF",  X"07",  X"07",  X"10",  X"10",  X"00",  X"10",  X"07",
  X"27",  X"BF",  X"07",  X"A5",  X"40",  X"BF",  X"0C",  X"10",
  X"10",  X"27",  X"BF",  X"10",  X"07",  X"10",  X"27",  X"27",
  X"00",  X"10",  X"07",  X"10",  X"BF",  X"07",  X"BF",  X"A5",
  X"A5",  X"BF",  X"10",  X"10",  X"10",  X"00",  X"10",  X"10",
  X"10",  X"00",  X"10",  X"A2",  X"BF",  X"07",  X"BF",  X"38",
  X"27",  X"27",  X"00",  X"10",  X"07",  X"10",  X"BF",  X"07",
  X"07",  X"A3",  X"80",  X"07",  X"00",  X"07",  X"BF",  X"27",
  X"A0",  X"80",  X"10",  X"10",  X"00",  X"10",  X"10",  X"00",
  X"10",  X"A2",  X"80",  X"07",  X"A0",  X"80",  X"00",  X"27",
  X"07",  X"2C",  X"BF",  X"04",  X"80",  X"4C",  X"07",  X"88",
  X"BF",  X"4C",  X"80",  X"A0",  X"10",  X"4C",  X"A0",  X"BF",
  X"04",  X"BF",  X"10",  X"00",  X"BF",  X"28",  X"05",  X"27",
  X"27",  X"00",  X"10",  X"07",  X"00",  X"00",  X"10",  X"02",
  X"02",  X"00",  X"2A",  X"10",  X"10",  X"00",  X"10",  X"07",
  X"BF",  X"10",  X"10",  X"07",  X"20",  X"BF",  X"27",  X"07",
  X"A1",  X"80",  X"07",  X"03",  X"2C",  X"BF",  X"04",  X"10",
  X"2C",  X"BF",  X"04",  X"A1",  X"BF",  X"07",  X"3B",  X"20",
  X"30",  X"01",  X"2C",  X"BF",  X"04",  X"BF",  X"07",  X"07",
  X"88",  X"BF",  X"2C",  X"BF",  X"07",  X"A5",  X"10",  X"40",
  X"BF",  X"08",  X"BF",  X"A6",  X"BF",  X"00",  X"E3",  X"A6",
  X"80",  X"10",  X"16",  X"88",  X"80",  X"00",  X"10",  X"00",
  X"A2",  X"80",  X"16",  X"02",  X"A0",  X"80",  X"00",  X"16",
  X"28",  X"38",  X"88",  X"80",  X"30",  X"06",  X"A4",  X"80",
  X"88",  X"06",  X"26",  X"24",  X"80",  X"10",  X"06",  X"A4",
  X"80",  X"26",  X"80",  X"88",  X"24",  X"A4",  X"80",  X"16",
  X"06",  X"06",  X"10",  X"C0",  X"10",  X"A2",  X"BF",  X"04",
  X"16",  X"10",  X"10",  X"88",  X"80",  X"36",  X"00",  X"06",
  X"80",  X"10",  X"30",  X"88",  X"80",  X"10",  X"C7",  X"E8",
  X"88",  X"BF",  X"10",  X"00",  X"06",  X"10",  X"C7",  X"E8",
  X"00",  X"06",  X"BF",  X"10",  X"00",  X"00",  X"BF",  X"16",
  X"00",  X"10",  X"00",  X"E8",  X"00",  X"10",  X"12",  X"13",
  X"00",  X"10",  X"00",  X"10",  X"00",  X"13",  X"FF",  X"10",
  X"00",  X"E3",  X"16",  X"88",  X"80",  X"00",  X"00",  X"06",
  X"C7",  X"E8",  X"10",  X"12",  X"13",  X"00",  X"10",  X"00",
  X"E3",  X"10",  X"00",  X"10",  X"00",  X"12",  X"FF",  X"E8",
  X"00",  X"E3",  X"16",  X"88",  X"80",  X"00",  X"00",  X"06",
  X"C7",  X"E8",  X"10",  X"12",  X"13",  X"00",  X"10",  X"00",
  X"E3",  X"FF",  X"10",  X"10",  X"00",  X"00",  X"EE",  X"00",
  X"E3",  X"10",  X"10",  X"26",  X"10",  X"10",  X"26",  X"10",
  X"10",  X"26",  X"26",  X"36",  X"36",  X"26",  X"26",  X"26",
  X"26",  X"26",  X"26",  X"10",  X"10",  X"26",  X"07",  X"00",
  X"10",  X"10",  X"00",  X"10",  X"10",  X"00",  X"06",  X"00",
  X"10",  X"C7",  X"E8",  X"E3",  X"10",  X"10",  X"26",  X"10",
  X"26",  X"10",  X"06",  X"26",  X"26",  X"06",  X"26",  X"10",
  X"10",  X"FF",  X"10",  X"06",  X"10",  X"10",  X"10",  X"FF",
  X"10",  X"06",  X"10",  X"FF",  X"E8",  X"00",  X"E3",  X"2E",
  X"2E",  X"24",  X"2C",  X"10",  X"04",  X"FF",  X"04",  X"92",
  X"80",  X"06",  X"26",  X"26",  X"26",  X"10",  X"00",  X"10",
  X"C7",  X"E8",  X"E3",  X"FF",  X"00",  X"10",  X"00",  X"04",
  X"A0",  X"80",  X"00",  X"04",  X"04",  X"80",  X"80",  X"04",
  X"80",  X"04",  X"80",  X"04",  X"54",  X"A0",  X"BF",  X"80",
  X"10",  X"34",  X"10",  X"34",  X"07",  X"00",  X"10",  X"10",
  X"00",  X"10",  X"10",  X"00",  X"04",  X"00",  X"10",  X"FF",
  X"00",  X"24",  X"24",  X"24",  X"24",  X"24",  X"24",  X"24",
  X"24",  X"24",  X"24",  X"C7",  X"E8",  X"04",  X"A2",  X"80",
  X"10",  X"BF",  X"10",  X"FF",  X"10",  X"BF",  X"04",  X"FF",
  X"10",  X"A2",  X"BF",  X"24",  X"FF",  X"10",  X"10",  X"BF",
  X"26",  X"E3",  X"FF",  X"10",  X"10",  X"14",  X"04",  X"00",
  X"0C",  X"04",  X"20",  X"0E",  X"06",  X"A6",  X"80",  X"10",
  X"FF",  X"10",  X"04",  X"00",  X"A2",  X"80",  X"10",  X"10",
  X"FF",  X"10",  X"C7",  X"E8",  X"FF",  X"20",  X"A2",  X"80",
  X"24",  X"04",  X"14",  X"10",  X"20",  X"10",  X"10",  X"00",
  X"20",  X"FF",  X"20",  X"C7",  X"E8",  X"10",  X"FF",  X"10",
  X"04",  X"22",  X"A0",  X"BF",  X"10",  X"00",  X"22",  X"10",
  X"10",  X"20",  X"BF",  X"20",  X"E3",  X"A6",  X"80",  X"00",
  X"FF",  X"10",  X"06",  X"00",  X"0B",  X"10",  X"00",  X"11",
  X"00",  X"01",  X"A2",  X"80",  X"0B",  X"20",  X"8B",  X"80",
  X"10",  X"06",  X"20",  X"00",  X"00",  X"01",  X"A2",  X"80",
  X"10",  X"00",  X"22",  X"10",  X"22",  X"00",  X"02",  X"8A",
  X"80",  X"10",  X"A3",  X"80",  X"00",  X"00",  X"00",  X"23",
  X"20",  X"10",  X"20",  X"A3",  X"80",  X"20",  X"A0",  X"80",
  X"30",  X"30",  X"A0",  X"80",  X"00",  X"30",  X"03",  X"2B",
  X"01",  X"03",  X"A0",  X"80",  X"00",  X"80",  X"01",  X"A3",
  X"80",  X"00",  X"00",  X"09",  X"A0",  X"BF",  X"00",  X"00",
  X"20",  X"20",  X"20",  X"20",  X"FF",  X"E8",  X"C7",  X"E8",
  X"00",  X"10",  X"12",  X"A3",  X"BF",  X"00",  X"23",  X"23",
  X"20",  X"20",  X"10",  X"20",  X"20",  X"FF",  X"E8",  X"28",
  X"01",  X"00",  X"20",  X"20",  X"01",  X"23",  X"20",  X"38",
  X"10",  X"28",  X"13",  X"21",  X"FF",  X"E8",  X"8B",  X"80",
  X"03",  X"06",  X"20",  X"00",  X"00",  X"00",  X"23",  X"20",
  X"21",  X"10",  X"20",  X"10",  X"00",  X"A0",  X"BF",  X"10",
  X"00",  X"FF",  X"10",  X"FF",  X"E8",  X"A0",  X"BF",  X"2B",
  X"A0",  X"80",  X"A0",  X"30",  X"03",  X"BF",  X"2B",  X"3B",
  X"10",  X"28",  X"13",  X"21",  X"BF",  X"10",  X"80",  X"A0",
  X"30",  X"03",  X"BF",  X"2B",  X"10",  X"BF",  X"10",  X"30",
  X"03",  X"BF",  X"2B",  X"E3",  X"06",  X"A0",  X"80",  X"10",
  X"16",  X"88",  X"80",  X"10",  X"06",  X"A0",  X"80",  X"10",
  X"88",  X"06",  X"10",  X"80",  X"10",  X"A4",  X"80",  X"10",
  X"A4",  X"80",  X"10",  X"10",  X"04",  X"C0",  X"04",  X"A2",
  X"80",  X"24",  X"06",  X"20",  X"A0",  X"80",  X"26",  X"04",
  X"A4",  X"BF",  X"10",  X"04",  X"04",  X"BF",  X"04",  X"10",
  X"C7",  X"E8",  X"10",  X"88",  X"15",  X"80",  X"10",  X"10",
  X"10",  X"10",  X"A4",  X"80",  X"04",  X"A5",  X"80",  X"10",
  X"A5",  X"80",  X"10",  X"10",  X"04",  X"04",  X"02",  X"A5",
  X"80",  X"04",  X"04",  X"A2",  X"80",  X"A5",  X"10",  X"00",
  X"10",  X"04",  X"00",  X"24",  X"FF",  X"10",  X"A2",  X"80",
  X"14",  X"A5",  X"80",  X"00",  X"06",  X"20",  X"A0",  X"BF",
  X"26",  X"24",  X"A4",  X"BF",  X"05",  X"04",  X"04",  X"10",
  X"BF",  X"04",  X"04",  X"A4",  X"80",  X"10",  X"10",  X"10",
  X"10",  X"00",  X"10",  X"04",  X"04",  X"20",  X"00",  X"24",
  X"24",  X"10",  X"10",  X"06",  X"20",  X"A4",  X"BF",  X"26",
  X"14",  X"24",  X"05",  X"A4",  X"80",  X"04",  X"28",  X"30",
  X"88",  X"80",  X"04",  X"A4",  X"BF",  X"10",  X"88",  X"BF",
  X"04",  X"04",  X"04",  X"05",  X"25",  X"04",  X"00",  X"10",
  X"92",  X"80",  X"00",  X"24",  X"24",  X"24",  X"24",  X"10",
  X"BF",  X"10",  X"04",  X"BF",  X"04",  X"A4",  X"04",  X"80",
  X"10",  X"04",  X"A2",  X"80",  X"04",  X"10",  X"00",  X"10",
  X"04",  X"00",  X"24",  X"FF",  X"10",  X"A2",  X"BF",  X"06",
  X"14",  X"10",  X"34",  X"C7",  X"E8",  X"04",  X"A4",  X"80",
  X"10",  X"04",  X"04",  X"C0",  X"10",  X"92",  X"BF",  X"14",
  X"BF",  X"10",  X"00",  X"10",  X"04",  X"04",  X"20",  X"00",
  X"24",  X"24",  X"10",  X"BF",  X"10",  X"A5",  X"80",  X"10",
  X"04",  X"04",  X"C0",  X"10",  X"92",  X"BF",  X"14",  X"A5",
  X"BF",  X"06",  X"FF",  X"10",  X"A2",  X"BF",  X"10",  X"BF",
  X"06",  X"00",  X"10",  X"04",  X"04",  X"20",  X"00",  X"24",
  X"24",  X"BF",  X"10",  X"10",  X"10",  X"00",  X"04",  X"A2",
  X"BF",  X"10",  X"02",  X"BF",  X"25",  X"10",  X"FF",  X"10",
  X"A2",  X"BF",  X"00",  X"14",  X"BF",  X"10",  X"05",  X"FF",
  X"04",  X"BF",  X"14",  X"E3",  X"FF",  X"10",  X"84",  X"80",
  X"10",  X"04",  X"84",  X"80",  X"04",  X"80",  X"04",  X"54",
  X"10",  X"A0",  X"80",  X"10",  X"C6",  X"00",  X"14",  X"16",
  X"88",  X"80",  X"04",  X"84",  X"80",  X"04",  X"04",  X"14",
  X"28",  X"A0",  X"BF",  X"84",  X"30",  X"88",  X"BF",  X"54",
  X"04",  X"00",  X"10",  X"54",  X"A0",  X"BF",  X"14",  X"00",
  X"10",  X"84",  X"BF",  X"04",  X"04",  X"A4",  X"BF",  X"04",
  X"FF",  X"00",  X"C7",  X"E8",  X"E3",  X"FF",  X"00",  X"86",
  X"80",  X"10",  X"04",  X"84",  X"80",  X"04",  X"80",  X"04",
  X"54",  X"A0",  X"80",  X"10",  X"C6",  X"00",  X"14",  X"16",
  X"88",  X"80",  X"04",  X"84",  X"80",  X"04",  X"04",  X"14",
  X"28",  X"A0",  X"BF",  X"84",  X"30",  X"88",  X"BF",  X"54",
  X"04",  X"00",  X"10",  X"54",  X"A0",  X"BF",  X"14",  X"00",
  X"10",  X"84",  X"BF",  X"04",  X"04",  X"A4",  X"BF",  X"04",
  X"FF",  X"00",  X"C7",  X"E8",  X"10",  X"C3",  X"00",  X"10",
  X"C3",  X"12",  X"10",  X"C3",  X"12",  X"E3",  X"10",  X"A6",
  X"10",  X"80",  X"16",  X"10",  X"10",  X"00",  X"10",  X"A2",
  X"80",  X"10",  X"24",  X"24",  X"C7",  X"EC",  X"10",  X"10",
  X"00",  X"12",  X"A2",  X"BF",  X"24",  X"C7",  X"E8",  X"10",
  X"10",  X"00",  X"10",  X"10",  X"13",  X"FF",  X"10",  X"00",
  X"E3",  X"16",  X"88",  X"80",  X"06",  X"56",  X"A2",  X"80",
  X"10",  X"04",  X"00",  X"07",  X"A2",  X"80",  X"17",  X"00",
  X"08",  X"00",  X"18",  X"A0",  X"00",  X"60",  X"A0",  X"80",
  X"06",  X"16",  X"10",  X"80",  X"36",  X"16",  X"10",  X"10",
  X"36",  X"04",  X"FF",  X"10",  X"A2",  X"80",  X"10",  X"16",
  X"00",  X"10",  X"26",  X"26",  X"36",  X"10",  X"10",  X"20",
  X"10",  X"A4",  X"80",  X"26",  X"00",  X"56",  X"A2",  X"80",
  X"00",  X"16",  X"10",  X"36",  X"C7",  X"E8",  X"26",  X"26",
  X"10",  X"26",  X"C7",  X"E8",  X"10",  X"10",  X"A0",  X"BF",
  X"16",  X"10",  X"10",  X"26",  X"BF",  X"36",  X"16",  X"10",
  X"06",  X"26",  X"26",  X"36",  X"10",  X"26",  X"C7",  X"E8",
  X"E3",  X"0E",  X"A6",  X"80",  X"10",  X"8E",  X"80",  X"2E",
  X"3F",  X"03",  X"20",  X"2B",  X"11",  X"03",  X"10",  X"2B",
  X"03",  X"06",  X"1B",  X"00",  X"28",  X"88",  X"80",  X"06",
  X"0E",  X"A0",  X"80",  X"00",  X"0E",  X"A0",  X"80",  X"06",
  X"0E",  X"A0",  X"80",  X"06",  X"0E",  X"A0",  X"80",  X"06",
  X"A6",  X"BF",  X"06",  X"10",  X"A6",  X"80",  X"08",  X"C7",
  X"E8",  X"A6",  X"BF",  X"00",  X"08",  X"A0",  X"BF",  X"06",
  X"C7",  X"E8",  X"C7",  X"E8",  X"E3",  X"A6",  X"10",  X"10",
  X"80",  X"10",  X"16",  X"88",  X"80",  X"10",  X"A0",  X"80",
  X"10",  X"09",  X"2B",  X"00",  X"A0",  X"BF",  X"09",  X"C7",
  X"E8",  X"10",  X"00",  X"20",  X"00",  X"A0",  X"00",  X"20",
  X"00",  X"20",  X"00",  X"20",  X"00",  X"BF",  X"00",  X"06",
  X"36",  X"2B",  X"03",  X"26",  X"2B",  X"A6",  X"06",  X"10",
  X"BF",  X"06",  X"10",  X"01",  X"23",  X"00",  X"26",  X"A0",
  X"BF",  X"01",  X"06",  X"36",  X"28",  X"00",  X"26",  X"28",
  X"01",  X"BF",  X"03",  X"E3",  X"A6",  X"10",  X"10",  X"80",
  X"10",  X"06",  X"A6",  X"80",  X"A6",  X"A6",  X"80",  X"06",
  X"06",  X"00",  X"08",  X"00",  X"00",  X"A0",  X"BF",  X"28",
  X"C7",  X"E8",  X"A6",  X"80",  X"16",  X"A0",  X"BF",  X"10",
  X"09",  X"2B",  X"00",  X"A0",  X"BF",  X"09",  X"C7",  X"E8",
  X"88",  X"BF",  X"A0",  X"10",  X"10",  X"10",  X"00",  X"20",
  X"00",  X"A0",  X"00",  X"20",  X"00",  X"20",  X"00",  X"20",
  X"00",  X"BF",  X"00",  X"06",  X"36",  X"2B",  X"03",  X"26",
  X"2B",  X"A6",  X"06",  X"10",  X"BF",  X"06",  X"10",  X"01",
  X"23",  X"00",  X"26",  X"A0",  X"BF",  X"01",  X"06",  X"36",
  X"28",  X"00",  X"26",  X"28",  X"01",  X"BF",  X"03",  X"E3",
  X"0E",  X"A6",  X"80",  X"10",  X"8E",  X"80",  X"10",  X"28",
  X"10",  X"A6",  X"28",  X"10",  X"10",  X"10",  X"80",  X"10",
  X"20",  X"20",  X"20",  X"20",  X"01",  X"A1",  X"BF",  X"00",
  X"06",  X"08",  X"08",  X"A6",  X"03",  X"80",  X"06",  X"10",
  X"23",  X"00",  X"26",  X"A1",  X"BF",  X"23",  X"06",  X"08",
  X"08",  X"00",  X"03",  X"10",  X"A6",  X"80",  X"10",  X"28",
  X"00",  X"A0",  X"BF",  X"28",  X"C7",  X"E8",  X"A2",  X"80",
  X"00",  X"02",  X"02",  X"28",  X"00",  X"22",  X"20",  X"C3",
  X"00",  X"10",  X"3F",  X"8A",  X"80",  X"10",  X"28",  X"10",
  X"3F",  X"88",  X"80",  X"3C",  X"02",  X"28",  X"88",  X"80",
  X"30",  X"02",  X"28",  X"88",  X"80",  X"A0",  X"02",  X"28",
  X"A0",  X"80",  X"10",  X"88",  X"80",  X"02",  X"C3",  X"00",
  X"C3",  X"10",  X"02",  X"88",  X"80",  X"00",  X"88",  X"80",
  X"10",  X"88",  X"80",  X"10",  X"30",  X"22",  X"C3",  X"10",
  X"10",  X"88",  X"80",  X"10",  X"88",  X"80",  X"88",  X"00",
  X"30",  X"88",  X"80",  X"88",  X"00",  X"30",  X"88",  X"80",
  X"88",  X"00",  X"30",  X"88",  X"80",  X"22",  X"30",  X"A0",
  X"80",  X"00",  X"22",  X"C3",  X"10",  X"30",  X"88",  X"BF",
  X"10",  X"BF",  X"00",  X"10",  X"C3",  X"10",  X"30",  X"10",
  X"22",  X"C3",  X"10",  X"E3",  X"10",  X"06",  X"06",  X"A6",
  X"80",  X"00",  X"28",  X"06",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"A3",  X"80",  X"A0",  X"BF",
  X"00",  X"C7",  X"E8",  X"A3",  X"60",  X"16",  X"C7",  X"E8",
  X"1F",  X"3F",  X"0A",  X"00",  X"A0",  X"80",  X"03",  X"10",
  X"10",  X"3B",  X"1B",  X"C3",  X"23",  X"20",  X"38",  X"A0",
  X"80",  X"00",  X"00",  X"A0",  X"80",  X"10",  X"10",  X"10",
  X"3B",  X"1B",  X"C3",  X"23",  X"38",  X"10",  X"29",  X"BF",
  X"10",  X"10",  X"39",  X"3B",  X"1B",  X"C3",  X"23",  X"E3",
  X"06",  X"04",  X"2C",  X"06",  X"FF",  X"10",  X"10",  X"20",
  X"26",  X"06",  X"A2",  X"80",  X"06",  X"10",  X"A6",  X"20",
  X"80",  X"10",  X"04",  X"30",  X"34",  X"02",  X"0F",  X"2C",
  X"13",  X"10",  X"3F",  X"1F",  X"C7",  X"E8",  X"A6",  X"80",
  X"10",  X"82",  X"80",  X"0F",  X"10",  X"A4",  X"20",  X"80",
  X"10",  X"04",  X"31",  X"28",  X"30",  X"0F",  X"2C",  X"11",
  X"12",  X"12",  X"3F",  X"1F",  X"C7",  X"E8",  X"0F",  X"10",
  X"14",  X"3F",  X"1F",  X"C7",  X"E8",  X"04",  X"82",  X"BF",
  X"04",  X"BF",  X"10",  X"E3",  X"07",  X"FF",  X"10",  X"A0",
  X"07",  X"10",  X"27",  X"FF",  X"27",  X"06",  X"06",  X"07",
  X"07",  X"21",  X"20",  X"07",  X"28",  X"07",  X"00",  X"A0",
  X"80",  X"A0",  X"27",  X"28",  X"07",  X"00",  X"27",  X"07",
  X"A0",  X"A2",  X"C7",  X"E8",  X"27",  X"28",  X"07",  X"20",
  X"27",  X"07",  X"A0",  X"A2",  X"C7",  X"E8",  X"A2",  X"80",
  X"10",  X"18",  X"10",  X"18",  X"82",  X"BF",  X"A0",  X"C3",
  X"00",  X"2A",  X"10",  X"10",  X"C3",  X"18",  X"E3",  X"06",
  X"A0",  X"80",  X"10",  X"2E",  X"00",  X"A6",  X"80",  X"10",
  X"06",  X"20",  X"26",  X"26",  X"C7",  X"E8",  X"10",  X"10",
  X"00",  X"10",  X"24",  X"10",  X"A2",  X"BF",  X"10",  X"C7",
  X"E8",  X"10",  X"10",  X"2C",  X"04",  X"00",  X"2A",  X"92",
  X"BF",  X"00",  X"26",  X"26",  X"26",  X"26",  X"C7",  X"E8",
  X"E3",  X"10",  X"10",  X"27",  X"FF",  X"27",  X"3F",  X"2E",
  X"27",  X"20",  X"10",  X"2E",  X"30",  X"A4",  X"80",  X"10",
  X"00",  X"10",  X"27",  X"A4",  X"80",  X"00",  X"27",  X"FF",
  X"07",  X"A2",  X"80",  X"07",  X"07",  X"26",  X"07",  X"A0",
  X"26",  X"40",  X"04",  X"A4",  X"80",  X"26",  X"02",  X"04",
  X"26",  X"28",  X"06",  X"FF",  X"00",  X"2C",  X"24",  X"27",
  X"C7",  X"E8",  X"FF",  X"07",  X"07",  X"26",  X"10",  X"26",
  X"02",  X"A4",  X"BF",  X"10",  X"04",  X"04",  X"26",  X"10",
  X"20",  X"27",  X"C7",  X"E8",  X"07",  X"20",  X"28",  X"10",
  X"26",  X"30",  X"BF",  X"27",  X"E3",  X"06",  X"06",  X"A4",
  X"80",  X"10",  X"A4",  X"80",  X"10",  X"10",  X"06",  X"FF",
  X"06",  X"06",  X"06",  X"01",  X"22",  X"28",  X"02",  X"06",
  X"2A",  X"00",  X"06",  X"06",  X"02",  X"13",  X"06",  X"02",
  X"10",  X"06",  X"04",  X"33",  X"0B",  X"30",  X"08",  X"22",
  X"20",  X"00",  X"38",  X"02",  X"30",  X"06",  X"30",  X"04",
  X"00",  X"A2",  X"BF",  X"38",  X"A4",  X"80",  X"00",  X"00",
  X"13",  X"04",  X"30",  X"08",  X"00",  X"38",  X"00",  X"30",
  X"04",  X"30",  X"A6",  X"00",  X"BF",  X"38",  X"00",  X"A0",
  X"80",  X"00",  X"00",  X"00",  X"A0",  X"BF",  X"01",  X"22",
  X"C7",  X"E8",  X"00",  X"06",  X"28",  X"06",  X"06",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"A1",  X"80",  X"A4",
  X"BF",  X"00",  X"FF",  X"10",  X"10",  X"22",  X"22",  X"C7",
  X"E8",  X"A1",  X"BF",  X"10",  X"10",  X"10",  X"10",  X"BF",
  X"06",  X"E3",  X"06",  X"06",  X"04",  X"3E",  X"10",  X"04",
  X"A4",  X"80",  X"06",  X"28",  X"A4",  X"BF",  X"02",  X"FF",
  X"10",  X"A4",  X"80",  X"02",  X"10",  X"20",  X"00",  X"A0",
  X"BF",  X"00",  X"00",  X"28",  X"02",  X"00",  X"06",  X"01",
  X"8E",  X"29",  X"06",  X"06",  X"80",  X"01",  X"10",  X"10",
  X"23",  X"00",  X"2B",  X"10",  X"20",  X"00",  X"00",  X"00",
  X"A1",  X"BF",  X"30",  X"20",  X"A0",  X"40",  X"04",  X"06",
  X"28",  X"00",  X"26",  X"04",  X"20",  X"22",  X"C7",  X"E8",
  X"00",  X"20",  X"00",  X"A1",  X"BF",  X"00",  X"00",  X"20",
  X"00",  X"A1",  X"BF",  X"00",  X"BF",  X"04",  X"E3",  X"06",
  X"06",  X"A4",  X"80",  X"10",  X"10",  X"10",  X"10",  X"06",
  X"04",  X"A5",  X"80",  X"06",  X"02",  X"FF",  X"05",  X"02",
  X"2D",  X"02",  X"05",  X"A6",  X"80",  X"10",  X"10",  X"20",
  X"00",  X"A5",  X"BF",  X"20",  X"04",  X"2D",  X"06",  X"06",
  X"27",  X"04",  X"06",  X"2F",  X"06",  X"07",  X"A7",  X"80",
  X"05",  X"00",  X"14",  X"07",  X"88",  X"80",  X"27",  X"07",
  X"10",  X"10",  X"06",  X"07",  X"00",  X"0D",  X"04",  X"07",
  X"0C",  X"02",  X"00",  X"35",  X"04",  X"34",  X"34",  X"02",
  X"04",  X"34",  X"06",  X"34",  X"A5",  X"04",  X"BF",  X"36",
  X"24",  X"07",  X"30",  X"A0",  X"80",  X"27",  X"06",  X"07",
  X"10",  X"10",  X"10",  X"06",  X"07",  X"0D",  X"00",  X"34",
  X"04",  X"04",  X"34",  X"07",  X"34",  X"35",  X"00",  X"34",
  X"04",  X"04",  X"06",  X"0C",  X"A5",  X"02",  X"06",  X"BF",
  X"36",  X"24",  X"07",  X"A7",  X"BF",  X"06",  X"A5",  X"80",
  X"26",  X"05",  X"A0",  X"80",  X"05",  X"26",  X"C7",  X"E8",
  X"05",  X"A0",  X"80",  X"26",  X"85",  X"BF",  X"05",  X"26",
  X"C7",  X"E8",  X"10",  X"10",  X"BF",  X"10",  X"E3",  X"10",
  X"FF",  X"10",  X"10",  X"22",  X"22",  X"C7",  X"E8",  X"E3",
  X"06",  X"00",  X"06",  X"15",  X"10",  X"04",  X"0D",  X"00",
  X"10",  X"35",  X"06",  X"00",  X"10",  X"34",  X"0C",  X"06",
  X"2E",  X"00",  X"24",  X"04",  X"04",  X"A4",  X"BF",  X"36",
  X"A6",  X"80",  X"00",  X"06",  X"A4",  X"80",  X"06",  X"04",
  X"28",  X"06",  X"04",  X"26",  X"20",  X"C7",  X"E8",  X"02",
  X"FF",  X"10",  X"06",  X"10",  X"06",  X"02",  X"02",  X"FF",
  X"2A",  X"06",  X"06",  X"28",  X"00",  X"26",  X"20",  X"BF",
  X"10",  X"E3",  X"8E",  X"80",  X"10",  X"3E",  X"A6",  X"80",
  X"00",  X"04",  X"A4",  X"80",  X"10",  X"8E",  X"80",  X"10",
  X"3E",  X"A6",  X"80",  X"00",  X"04",  X"A2",  X"80",  X"10",
  X"10",  X"8E",  X"BF",  X"3E",  X"10",  X"10",  X"FF",  X"10",
  X"A6",  X"80",  X"3E",  X"04",  X"06",  X"28",  X"00",  X"26",
  X"20",  X"A6",  X"BF",  X"10",  X"C7",  X"E8",  X"10",  X"FF",
  X"10",  X"24",  X"22",  X"BF",  X"10",  X"00",  X"10",  X"28",
  X"10",  X"00",  X"10",  X"10",  X"FF",  X"10",  X"BF",  X"10",
  X"FF",  X"10",  X"24",  X"10",  X"BF",  X"22",  X"E3",  X"10",
  X"00",  X"06",  X"10",  X"A2",  X"10",  X"80",  X"10",  X"28",
  X"A2",  X"BF",  X"02",  X"FF",  X"10",  X"10",  X"22",  X"22",
  X"A6",  X"06",  X"80",  X"10",  X"06",  X"4E",  X"10",  X"02",
  X"10",  X"FF",  X"10",  X"04",  X"A6",  X"BF",  X"4E",  X"04",
  X"10",  X"04",  X"A6",  X"80",  X"10",  X"4C",  X"10",  X"02",
  X"10",  X"FF",  X"10",  X"06",  X"06",  X"A6",  X"BF",  X"4C",
  X"C7",  X"E8",  X"E3",  X"A6",  X"80",  X"10",  X"FF",  X"E8",
  X"FF",  X"10",  X"06",  X"05",  X"06",  X"A4",  X"80",  X"10",
  X"10",  X"10",  X"A4",  X"80",  X"10",  X"C7",  X"E8",  X"0C",
  X"10",  X"A4",  X"BF",  X"34",  X"89",  X"BF",  X"08",  X"A5",
  X"80",  X"10",  X"10",  X"15",  X"05",  X"05",  X"A1",  X"80",
  X"04",  X"00",  X"0D",  X"00",  X"03",  X"8B",  X"80",  X"10",
  X"0D",  X"05",  X"A4",  X"80",  X"00",  X"88",  X"80",  X"A0",
  X"06",  X"25",  X"04",  X"80",  X"0C",  X"A0",  X"80",  X"04",
  X"05",  X"A4",  X"80",  X"00",  X"10",  X"A4",  X"80",  X"10",
  X"04",  X"04",  X"05",  X"04",  X"20",  X"A2",  X"80",  X"20",
  X"A2",  X"10",  X"80",  X"10",  X"06",  X"24",  X"A2",  X"04",
  X"06",  X"24",  X"80",  X"06",  X"06",  X"24",  X"A2",  X"04",
  X"00",  X"24",  X"80",  X"00",  X"00",  X"24",  X"04",  X"00",
  X"24",  X"00",  X"00",  X"20",  X"10",  X"10",  X"00",  X"20",
  X"00",  X"20",  X"80",  X"04",  X"10",  X"05",  X"24",  X"A0",
  X"80",  X"00",  X"08",  X"10",  X"20",  X"00",  X"04",  X"10",
  X"24",  X"FF",  X"10",  X"C7",  X"E8",  X"08",  X"10",  X"20",
  X"10",  X"22",  X"02",  X"10",  X"00",  X"10",  X"20",  X"FF",
  X"02",  X"BF",  X"BF",  X"10",  X"00",  X"05",  X"10",  X"21",
  X"10",  X"BF",  X"20",  X"04",  X"04",  X"05",  X"A5",  X"BF",
  X"A4",  X"04",  X"04",  X"05",  X"04",  X"20",  X"A2",  X"80",
  X"20",  X"A2",  X"10",  X"80",  X"10",  X"06",  X"24",  X"A2",
  X"04",  X"06",  X"24",  X"80",  X"06",  X"06",  X"24",  X"A2",
  X"04",  X"00",  X"24",  X"80",  X"00",  X"00",  X"24",  X"04",
  X"00",  X"24",  X"00",  X"00",  X"20",  X"00",  X"20",  X"00",
  X"20",  X"04",  X"25",  X"10",  X"20",  X"25",  X"10",  X"04",
  X"08",  X"14",  X"FF",  X"24",  X"C7",  X"E8",  X"10",  X"FF",
  X"10",  X"92",  X"80",  X"06",  X"05",  X"08",  X"05",  X"A0",
  X"80",  X"05",  X"A2",  X"80",  X"A2",  X"10",  X"80",  X"10",
  X"06",  X"26",  X"A2",  X"06",  X"06",  X"26",  X"80",  X"06",
  X"06",  X"26",  X"A2",  X"06",  X"06",  X"26",  X"80",  X"06",
  X"06",  X"26",  X"06",  X"06",  X"06",  X"26",  X"00",  X"20",
  X"00",  X"20",  X"00",  X"20",  X"10",  X"FF",  X"10",  X"FF",
  X"10",  X"C7",  X"E8",  X"00",  X"05",  X"04",  X"20",  X"20",
  X"A2",  X"04",  X"04",  X"20",  X"BF",  X"20",  X"10",  X"FF",
  X"10",  X"10",  X"BF",  X"04",  X"01",  X"0D",  X"05",  X"A3",
  X"BF",  X"10",  X"05",  X"23",  X"10",  X"20",  X"25",  X"10",
  X"05",  X"08",  X"14",  X"FF",  X"25",  X"C7",  X"E8",  X"FF",
  X"10",  X"BF",  X"10",  X"BF",  X"04",  X"00",  X"0C",  X"10",
  X"04",  X"BF",  X"05",  X"10",  X"FF",  X"10",  X"BF",  X"04",
  X"E3",  X"A6",  X"80",  X"10",  X"06",  X"A4",  X"80",  X"06",
  X"04",  X"80",  X"80",  X"04",  X"00",  X"2C",  X"04",  X"04",
  X"C0",  X"04",  X"84",  X"BF",  X"04",  X"04",  X"A4",  X"BF",
  X"04",  X"06",  X"A0",  X"80",  X"00",  X"C0",  X"10",  X"C7",
  X"E8",  X"BF",  X"00",  X"E3",  X"06",  X"A2",  X"80",  X"00",
  X"FF",  X"10",  X"FF",  X"E8",  X"00",  X"E3",  X"10",  X"00",
  X"A6",  X"80",  X"00",  X"06",  X"A2",  X"80",  X"06",  X"10",
  X"02",  X"A4",  X"80",  X"04",  X"10",  X"10",  X"FF",  X"04",
  X"A4",  X"BF",  X"10",  X"06",  X"04",  X"A4",  X"BF",  X"02",
  X"FF",  X"10",  X"06",  X"A4",  X"80",  X"06",  X"06",  X"A4",
  X"80",  X"06",  X"10",  X"10",  X"FF",  X"04",  X"A4",  X"BF",
  X"10",  X"06",  X"A2",  X"80",  X"06",  X"FF",  X"10",  X"06",
  X"A0",  X"80",  X"06",  X"C7",  X"E8",  X"C0",  X"10",  X"06",
  X"A6",  X"BF",  X"00",  X"FF",  X"E8",  X"00",  X"20",  X"1F",
  X"10",  X"20",  X"30",  X"2A",  X"10",  X"20",  X"20",  X"12",
  X"38",  X"C3",  X"02",  X"20",  X"2A",  X"20",  X"12",  X"32",
  X"12",  X"1F",  X"20",  X"C3",  X"32",  X"52",  X"10",  X"00",
  X"13",  X"00",  X"10",  X"00",  X"E3",  X"10",  X"56",  X"00",
  X"10",  X"00",  X"10",  X"A2",  X"80",  X"00",  X"16",  X"10",
  X"26",  X"36",  X"C7",  X"E8",  X"16",  X"00",  X"28",  X"36",
  X"C7",  X"E8",  X"E3",  X"16",  X"10",  X"88",  X"10",  X"10",
  X"80",  X"10",  X"04",  X"56",  X"10",  X"00",  X"10",  X"16",
  X"00",  X"28",  X"04",  X"54",  X"34",  X"00",  X"E8",  X"00",
  X"E3",  X"10",  X"56",  X"00",  X"10",  X"00",  X"10",  X"A2",
  X"80",  X"16",  X"06",  X"00",  X"26",  X"C7",  X"E8",  X"00",
  X"28",  X"36",  X"C7",  X"E8",  X"12",  X"88",  X"80",  X"4A",
  X"02",  X"02",  X"A0",  X"80",  X"3F",  X"20",  X"10",  X"10",
  X"10",  X"00",  X"28",  X"88",  X"80",  X"02",  X"C3",  X"10",
  X"28",  X"88",  X"80",  X"10",  X"02",  X"02",  X"02",  X"02",
  X"A0",  X"BF",  X"00",  X"4A",  X"A0",  X"80",  X"0A",  X"80",
  X"0A",  X"02",  X"4A",  X"02",  X"A0",  X"80",  X"0A",  X"4A",
  X"A0",  X"BF",  X"0A",  X"08",  X"08",  X"C3",  X"20",  X"0A",
  X"08",  X"08",  X"C3",  X"20",  X"C3",  X"00",  X"E3",  X"8E",
  X"80",  X"10",  X"06",  X"3F",  X"13",  X"00",  X"28",  X"20",
  X"11",  X"88",  X"80",  X"10",  X"00",  X"00",  X"00",  X"28",
  X"88",  X"80",  X"48",  X"00",  X"00",  X"00",  X"28",  X"88",
  X"BF",  X"00",  X"80",  X"48",  X"48",  X"A0",  X"BF",  X"00",
  X"20",  X"C7",  X"E8",  X"E3",  X"10",  X"10",  X"10",  X"24",
  X"00",  X"10",  X"A2",  X"80",  X"04",  X"C7",  X"E8",  X"A0",
  X"BF",  X"00",  X"26",  X"C7",  X"E8",  X"E3",  X"10",  X"00",
  X"10",  X"10",  X"FF",  X"10",  X"92",  X"80",  X"00",  X"06",
  X"0A",  X"02",  X"A2",  X"80",  X"A2",  X"80",  X"10",  X"26",
  X"26",  X"A2",  X"80",  X"06",  X"26",  X"26",  X"A2",  X"80",
  X"06",  X"26",  X"26",  X"06",  X"20",  X"20",  X"20",  X"C7",
  X"E8",  X"FF",  X"10",  X"C7",  X"E8",  X"E3",  X"10",  X"10",
  X"00",  X"24",  X"A2",  X"80",  X"04",  X"C7",  X"E8",  X"A0",
  X"BF",  X"00",  X"26",  X"C7",  X"E8",  X"E3",  X"A6",  X"80",
  X"10",  X"FF",  X"06",  X"16",  X"88",  X"80",  X"00",  X"10",
  X"04",  X"A2",  X"80",  X"16",  X"02",  X"A0",  X"80",  X"00",
  X"16",  X"28",  X"A0",  X"80",  X"30",  X"88",  X"80",  X"10",
  X"06",  X"A0",  X"80",  X"16",  X"C0",  X"06",  X"A2",  X"80",
  X"10",  X"16",  X"88",  X"80",  X"06",  X"06",  X"A2",  X"80",
  X"06",  X"A2",  X"80",  X"26",  X"FF",  X"04",  X"26",  X"06",
  X"A2",  X"80",  X"36",  X"FF",  X"04",  X"26",  X"36",  X"00",
  X"10",  X"00",  X"10",  X"FF",  X"00",  X"C7",  X"E8",  X"00",
  X"10",  X"BF",  X"10",  X"00",  X"10",  X"FF",  X"10",  X"C7",
  X"E8",  X"FF",  X"00",  X"16",  X"28",  X"A0",  X"BF",  X"30",
  X"BF",  X"FF",  X"10",  X"BF",  X"06",  X"FF",  X"10",  X"BF",
  X"10",  X"10",  X"10",  X"00",  X"13",  X"FF",  X"10",  X"00",
  X"E3",  X"10",  X"10",  X"10",  X"00",  X"24",  X"A2",  X"80",
  X"04",  X"C7",  X"E8",  X"A0",  X"BF",  X"00",  X"26",  X"C7",
  X"E8",  X"E3",  X"10",  X"10",  X"10",  X"24",  X"00",  X"10",
  X"A2",  X"80",  X"04",  X"C7",  X"E8",  X"A0",  X"BF",  X"00",
  X"26",  X"C7",  X"E8",  X"E3",  X"10",  X"10",  X"10",  X"24",
  X"00",  X"10",  X"A2",  X"80",  X"04",  X"C7",  X"E8",  X"A0",
  X"BF",  X"00",  X"26",  X"C7",  X"E8",  X"12",  X"82",  X"AB",
  X"80",  X"88",  X"23",  X"23",  X"23",  X"23",  X"23",  X"23",
  X"23",  X"23",  X"23",  X"23",  X"23",  X"23",  X"23",  X"23",
  X"23",  X"23",  X"23",  X"23",  X"23",  X"23",  X"23",  X"23",
  X"23",  X"23",  X"23",  X"23",  X"23",  X"23",  X"23",  X"23",
  X"23",  X"23",  X"23",  X"C3",  X"40",  X"23",  X"23",  X"23",
  X"23",  X"23",  X"23",  X"23",  X"23",  X"23",  X"23",  X"23",
  X"23",  X"23",  X"40",  X"2B",  X"33",  X"C3",  X"13",  X"80",
  X"10",  X"92",  X"80",  X"1A",  X"92",  X"80",  X"92",  X"80",
  X"20",  X"20",  X"92",  X"80",  X"10",  X"D0",  X"C3",  X"10",
  X"A2",  X"80",  X"10",  X"02",  X"A2",  X"80",  X"10",  X"A3",
  X"80",  X"10",  X"2B",  X"BF",  X"03",  X"83",  X"80",  X"00",
  X"28",  X"33",  X"03",  X"80",  X"20",  X"A3",  X"BF",  X"00",
  X"80",  X"00",  X"A0",  X"80",  X"00",  X"22",  X"10",  X"80",
  X"00",  X"2A",  X"80",  X"33",  X"22",  X"80",  X"02",  X"02",
  X"22",  X"A0",  X"BF",  X"92",  X"80",  X"2B",  X"A3",  X"BF",
  X"83",  X"80",  X"23",  X"92",  X"2A",  X"80",  X"33",  X"A2",
  X"80",  X"33",  X"A2",  X"80",  X"33",  X"A2",  X"80",  X"33",
  X"A2",  X"80",  X"02",  X"82",  X"80",  X"02",  X"82",  X"80",
  X"33",  X"A2",  X"80",  X"02",  X"82",  X"80",  X"02",  X"82",
  X"80",  X"33",  X"A2",  X"80",  X"33",  X"A2",  X"80",  X"02",
  X"82",  X"80",  X"02",  X"82",  X"80",  X"33",  X"A2",  X"80",
  X"02",  X"82",  X"80",  X"02",  X"82",  X"80",  X"33",  X"A2",
  X"80",  X"33",  X"A2",  X"80",  X"33",  X"A2",  X"80",  X"02",
  X"82",  X"80",  X"02",  X"82",  X"80",  X"33",  X"A2",  X"80",
  X"02",  X"82",  X"80",  X"02",  X"82",  X"80",  X"33",  X"A2",
  X"80",  X"33",  X"A2",  X"80",  X"02",  X"82",  X"80",  X"02",
  X"82",  X"80",  X"33",  X"A2",  X"80",  X"02",  X"82",  X"80",
  X"02",  X"A3",  X"BF",  X"92",  X"80",  X"22",  X"90",  X"80",
  X"20",  X"C3",  X"10",  X"80",  X"10",  X"92",  X"80",  X"10",
  X"92",  X"80",  X"92",  X"80",  X"20",  X"20",  X"92",  X"80",
  X"10",  X"D0",  X"C3",  X"10",  X"A2",  X"80",  X"10",  X"02",
  X"A2",  X"80",  X"10",  X"A3",  X"80",  X"10",  X"2B",  X"BF",
  X"03",  X"83",  X"80",  X"00",  X"28",  X"33",  X"03",  X"80",
  X"20",  X"A3",  X"BF",  X"00",  X"80",  X"00",  X"A0",  X"80",
  X"00",  X"22",  X"10",  X"80",  X"00",  X"2A",  X"80",  X"33",
  X"22",  X"80",  X"02",  X"02",  X"22",  X"A0",  X"BF",  X"92",
  X"80",  X"2B",  X"A3",  X"BF",  X"83",  X"80",  X"23",  X"92",
  X"2A",  X"80",  X"33",  X"A2",  X"80",  X"33",  X"A2",  X"80",
  X"33",  X"A2",  X"80",  X"33",  X"A2",  X"80",  X"02",  X"82",
  X"80",  X"02",  X"82",  X"80",  X"33",  X"A2",  X"80",  X"02",
  X"82",  X"80",  X"02",  X"82",  X"80",  X"33",  X"A2",  X"80",
  X"33",  X"A2",  X"80",  X"02",  X"82",  X"80",  X"02",  X"82",
  X"80",  X"33",  X"A2",  X"80",  X"02",  X"82",  X"80",  X"02",
  X"82",  X"80",  X"33",  X"A2",  X"80",  X"33",  X"A2",  X"80",
  X"33",  X"A2",  X"80",  X"02",  X"82",  X"80",  X"02",  X"82",
  X"80",  X"33",  X"A2",  X"80",  X"02",  X"82",  X"80",  X"02",
  X"82",  X"80",  X"33",  X"A2",  X"80",  X"33",  X"A2",  X"80",
  X"02",  X"82",  X"80",  X"02",  X"82",  X"80",  X"33",  X"A2",
  X"80",  X"02",  X"82",  X"80",  X"02",  X"A3",  X"BF",  X"92",
  X"80",  X"02",  X"90",  X"80",  X"20",  X"C3",  X"10",  X"C3",
  X"10",  X"00",  X"10",  X"32",  X"C3",  X"22",  X"C3",  X"10",
  X"E3",  X"00",  X"10",  X"10",  X"22",  X"C7",  X"E8",  X"E3",
  X"A6",  X"80",  X"10",  X"80",  X"80",  X"00",  X"06",  X"A6",
  X"80",  X"00",  X"00",  X"00",  X"2E",  X"2A",  X"3A",  X"A2",
  X"BF",  X"A2",  X"C7",  X"EE",  X"C7",  X"E8",  X"10",  X"00",
  X"A0",  X"80",  X"10",  X"00",  X"20",  X"C3",  X"10",  X"10",
  X"00",  X"20",  X"20",  X"C3",  X"10",  X"E3",  X"A6",  X"80",
  X"10",  X"80",  X"0E",  X"00",  X"3A",  X"04",  X"A6",  X"80",
  X"00",  X"0E",  X"2A",  X"3A",  X"A0",  X"BF",  X"00",  X"00",
  X"10",  X"0E",  X"2A",  X"00",  X"3A",  X"04",  X"A6",  X"BF",
  X"0E",  X"C7",  X"E8",  X"10",  X"00",  X"00",  X"00",  X"88",
  X"BF",  X"0A",  X"20",  X"A2",  X"80",  X"00",  X"C3",  X"00",
  X"00",  X"88",  X"BF",  X"10",  X"20",  X"C3",  X"00",  X"10",
  X"00",  X"A0",  X"00",  X"80",  X"10",  X"00",  X"88",  X"BF",
  X"00",  X"00",  X"C3",  X"00",  X"50",  X"10",  X"34",  X"10",
  X"05",  X"2C",  X"15",  X"E0",  X"90",  X"00",  X"00",  X"00",
  X"3B",  X"3B",  X"3B",  X"3B",  X"3B",  X"3B",  X"3B",  X"3B",
  X"E8",  X"10",  X"C4",  X"CC",  X"00",  X"00",  X"00",  X"50",
  X"2C",  X"10",  X"05",  X"34",  X"15",  X"95",  X"00",  X"00",
  X"00",  X"E8",  X"E8",  X"1B",  X"1B",  X"1B",  X"1B",  X"1B",
  X"1B",  X"1B",  X"1B",  X"E0",  X"E0",  X"C4",  X"CC",  X"50",
  X"10",  X"C5",  X"00",  X"10",  X"14",  X"24",  X"8C",  X"00",
  X"00",  X"00",  X"E3",  X"E3",  X"E3",  X"E3",  X"E3",  X"E3",
  X"E3",  X"E8",  X"E8",  X"E8",  X"E8",  X"E8",  X"E8",  X"E8",
  X"10",  X"14",  X"24",  X"03",  X"04",  X"23",  X"23",  X"80",
  X"10",  X"10",  X"15",  X"25",  X"25",  X"25",  X"25",  X"25",
  X"25",  X"E8",  X"48",  X"10",  X"88",  X"00",  X"00",  X"00",
  X"10",  X"01",  X"E0",  X"21",  X"A9",  X"80",  X"00",  X"00",
  X"A1",  X"BF",  X"00",  X"10",  X"01",  X"E8",  X"A9",  X"80",
  X"00",  X"00",  X"21",  X"A1",  X"BF",  X"00",  X"E0",  X"10",
  X"15",  X"05",  X"05",  X"05",  X"05",  X"05",  X"25",  X"8C",
  X"00",  X"00",  X"00",  X"C4",  X"CC",  X"14",  X"8C",  X"00",
  X"00",  X"00",  X"C4",  X"CC",  X"A6",  X"80",  X"14",  X"8D",
  X"14",  X"80",  X"A6",  X"80",  X"0E",  X"2C",  X"15",  X"8D",
  X"80",  X"A6",  X"80",  X"48",  X"15",  X"8D",  X"00",  X"00",
  X"00",  X"80",  X"A6",  X"80",  X"48",  X"2D",  X"8D",  X"00",
  X"00",  X"00",  X"80",  X"A6",  X"80",  X"00",  X"BF",  X"D0",
  X"C4",  X"CC",  X"10",  X"C3",  X"D0",  X"10",  X"C3",  X"D0",
  X"10",  X"C3",  X"D0",  X"00",  X"14",  X"14",  X"8C",  X"00",
  X"00",  X"00",  X"48",  X"00",  X"8C",  X"80",  X"00",  X"D0",
  X"10",  X"15",  X"05",  X"10",  X"15",  X"05",  X"A5",  X"80",
  X"00",  X"A0",  X"80",  X"00",  X"3D",  X"3D",  X"3D",  X"3D",
  X"3D",  X"3D",  X"3D",  X"3D",  X"3D",  X"3D",  X"3D",  X"3D",
  X"3D",  X"3D",  X"3D",  X"3D",  X"2D",  X"10",  X"15",  X"25",
  X"A0",  X"80",  X"00",  X"1D",  X"1D",  X"1D",  X"1D",  X"1D",
  X"1D",  X"1D",  X"1D",  X"1D",  X"1D",  X"1D",  X"1D",  X"1D",
  X"1D",  X"1D",  X"1D",  X"0D",  X"8C",  X"00",  X"00",  X"00",
  X"C4",  X"CC",  X"C3",  X"00",  X"C3",  X"00",  X"C3",  X"00",
  X"25",  X"50",  X"10",  X"15",  X"10",  X"C5",  X"00",  X"10",
  X"12",  X"02",  X"02",  X"22",  X"2D",  X"2C",  X"12",  X"10",
  X"12",  X"02",  X"A0",  X"80",  X"12",  X"8A",  X"00",  X"00",
  X"00",  X"10",  X"00",  X"03",  X"14",  X"8A",  X"00",  X"00",
  X"00",  X"10",  X"12",  X"02",  X"22",  X"22",  X"80",  X"10",
  X"E3",  X"10",  X"2E",  X"13",  X"A6",  X"10",  X"80",  X"03",
  X"2E",  X"10",  X"A0",  X"13",  X"80",  X"06",  X"A0",  X"80",
  X"10",  X"80",  X"06",  X"80",  X"06",  X"00",  X"A0",  X"BF",
  X"A0",  X"23",  X"26",  X"20",  X"10",  X"C7",  X"E8",  X"26",
  X"C7",  X"E8",  X"2A",  X"10",  X"10",  X"00",  X"22",  X"C3",
  X"20",  X"E3",  X"10",  X"10",  X"00",  X"A0",  X"80",  X"00",
  X"A6",  X"80",  X"10",  X"2E",  X"10",  X"10",  X"00",  X"A4",
  X"80",  X"10",  X"10",  X"10",  X"10",  X"15",  X"15",  X"15",
  X"80",  X"14",  X"10",  X"00",  X"24",  X"05",  X"A0",  X"80",
  X"04",  X"C0",  X"00",  X"04",  X"04",  X"10",  X"C0",  X"10",
  X"05",  X"A0",  X"80",  X"04",  X"C0",  X"00",  X"04",  X"00",
  X"24",  X"04",  X"A4",  X"80",  X"00",  X"04",  X"A0",  X"BF",
  X"04",  X"05",  X"A0",  X"BF",  X"04",  X"A0",  X"BF",  X"10",
  X"04",  X"A4",  X"BF",  X"04",  X"C7",  X"E8",  X"00",  X"BF",
  X"0E",  X"10",  X"48",  X"34",  X"09",  X"A1",  X"80",  X"10",
  X"11",  X"20",  X"11",  X"21",  X"10",  X"11",  X"20",  X"11",
  X"21",  X"80",  X"10",  X"10",  X"00",  X"00",  X"A0",  X"80",
  X"00",  X"02",  X"3F",  X"08",  X"00",  X"10",  X"10",  X"10",
  X"10",  X"00",  X"00",  X"A0",  X"80",  X"00",  X"00",  X"10",
  X"10",  X"11",  X"21",  X"10",  X"10",  X"10",  X"00",  X"00",
  X"A0",  X"80",  X"00",  X"00",  X"10",  X"02",  X"10",  X"11",
  X"21",  X"10",  X"10",  X"10",  X"00",  X"00",  X"A0",  X"80",
  X"00",  X"00",  X"10",  X"10",  X"11",  X"21",  X"02",  X"32",
  X"0A",  X"21",  X"10",  X"C3",  X"00",  X"10",  X"10",  X"10",
  X"D0",  X"C3",  X"00",  X"E3",  X"10",  X"00",  X"10",  X"A0",
  X"80",  X"10",  X"10",  X"C0",  X"10",  X"10",  X"C7",  X"E8",
  X"E3",  X"10",  X"00",  X"A0",  X"80",  X"10",  X"C0",  X"10",
  X"10",  X"C7",  X"E8",  X"E3",  X"10",  X"00",  X"A0",  X"80",
  X"10",  X"C0",  X"10",  X"10",  X"C7",  X"E8",  X"E3",  X"10",
  X"00",  X"A0",  X"80",  X"10",  X"C0",  X"10",  X"10",  X"C7",
  X"E8",  X"E3",  X"10",  X"00",  X"A0",  X"80",  X"10",  X"C0",
  X"10",  X"10",  X"C7",  X"E8",  X"E3",  X"10",  X"00",  X"A0",
  X"80",  X"10",  X"C0",  X"10",  X"10",  X"C7",  X"E8",  X"E3",
  X"10",  X"00",  X"A0",  X"80",  X"10",  X"C0",  X"10",  X"10",
  X"C7",  X"E8",  X"E3",  X"10",  X"00",  X"10",  X"A0",  X"80",
  X"10",  X"10",  X"C0",  X"10",  X"10",  X"C7",  X"E8",  X"00",
  X"10",  X"10",  X"C0",  X"00",  X"10",  X"10",  X"98",  X"10",
  X"10",  X"C0",  X"00",  X"10",  X"10",  X"C0",  X"00",  X"48",
  X"31",  X"09",  X"A1",  X"80",  X"00",  X"44",  X"31",  X"A1",
  X"80",  X"00",  X"FF",  X"00",  X"FF",  X"00",  X"23",  X"FF",
  X"00",  X"10",  X"D0",  X"00",  X"00",  X"8C",  X"80",  X"2C",
  X"D0",  X"8C",  X"00",  X"00",  X"00",  X"C4",  X"CC",  X"C3",
  X"00",  X"C1",  X"00",  X"48",  X"34",  X"09",  X"A1",  X"80",
  X"00",  X"10",  X"14",  X"10",  X"24",  X"44",  X"80",  X"10",
  X"14",  X"10",  X"24",  X"20",  X"04",  X"34",  X"09",  X"10",
  X"14",  X"24",  X"01",  X"10",  X"14",  X"24",  X"10",  X"14",
  X"21",  X"24",  X"C3",  X"00",  X"C3",  X"00",  X"D0",  X"00",
  X"00",  X"00",  X"C4",  X"CC",  X"48",  X"30",  X"08",  X"A0",
  X"80",  X"00",  X"44",  X"00",  X"28",  X"80",  X"10",  X"10",
  X"C1",  X"00",  X"E3",  X"10",  X"10",  X"14",  X"14",  X"A4",
  X"80",  X"00",  X"04",  X"A2",  X"80",  X"04",  X"C2",  X"00",
  X"A4",  X"BF",  X"04",  X"C7",  X"E8",  X"27",  X"25",  X"25",
  X"25",  X"25",  X"3D",  X"3D",  X"3D",  X"40",  X"25",  X"3D",
  X"3D",  X"3D",  X"3D",  X"10",  X"00",  X"25",  X"05",  X"20",
  X"10",  X"2D",  X"8D",  X"80",  X"00",  X"34",  X"10",  X"00",
  X"2C",  X"14",  X"08",  X"E0",  X"90",  X"3B",  X"3B",  X"3B",
  X"3B",  X"3B",  X"3B",  X"3B",  X"3B",  X"E8",  X"C5",  X"10",
  X"10",  X"10",  X"00",  X"A0",  X"80",  X"00",  X"C0",  X"03",
  X"03",  X"10",  X"20",  X"8C",  X"10",  X"28",  X"10",  X"00",
  X"30",  X"10",  X"50",  X"88",  X"80",  X"28",  X"10",  X"00",
  X"30",  X"10",  X"08",  X"90",  X"03",  X"80",  X"1B",  X"1B",
  X"1B",  X"1B",  X"03",  X"1B",  X"1B",  X"1B",  X"03",  X"03",
  X"03",  X"E8",  X"1B",  X"1B",  X"1B",  X"1B",  X"1B",  X"1B",
  X"1B",  X"1B",  X"80",  X"E0",  X"03",  X"80",  X"1B",  X"1B",
  X"1B",  X"1B",  X"03",  X"1B",  X"1B",  X"1B",  X"03",  X"03",
  X"03",  X"8C",  X"00",  X"00",  X"00",  X"C4",  X"CC",  X"27",
  X"25",  X"00",  X"2C",  X"25",  X"3D",  X"3D",  X"3D",  X"40",
  X"25",  X"10",  X"00",  X"25",  X"05",  X"20",  X"20",  X"10",
  X"2D",  X"8D",  X"80",  X"00",  X"34",  X"10",  X"00",  X"2C",
  X"14",  X"08",  X"E0",  X"90",  X"3B",  X"3B",  X"3B",  X"3B",
  X"3B",  X"3B",  X"3B",  X"3B",  X"E8",  X"C5",  X"10",  X"10",
  X"10",  X"00",  X"A0",  X"80",  X"00",  X"C0",  X"03",  X"03",
  X"10",  X"20",  X"10",  X"00",  X"A0",  X"80",  X"00",  X"03",
  X"00",  X"08",  X"2C",  X"14",  X"80",  X"03",  X"A0",  X"80",
  X"10",  X"20",  X"8C",  X"10",  X"28",  X"10",  X"00",  X"30",
  X"10",  X"50",  X"88",  X"80",  X"28",  X"10",  X"00",  X"30",
  X"10",  X"08",  X"90",  X"03",  X"80",  X"03",  X"1B",  X"1B",
  X"1B",  X"E8",  X"1B",  X"1B",  X"1B",  X"1B",  X"1B",  X"1B",
  X"1B",  X"1B",  X"80",  X"E0",  X"03",  X"80",  X"03",  X"1B",
  X"1B",  X"1B",  X"8C",  X"00",  X"00",  X"00",  X"C4",  X"CC",
  X"10",  X"10",  X"10",  X"2A",  X"03",  X"03",  X"32",  X"A2",
  X"80",  X"02",  X"32",  X"0A",  X"A2",  X"80",  X"10",  X"02",
  X"A2",  X"BF",  X"2A",  X"10",  X"C3",  X"10",  X"10",  X"10",
  X"2B",  X"00",  X"00",  X"32",  X"A2",  X"80",  X"03",  X"32",
  X"0A",  X"A2",  X"80",  X"10",  X"03",  X"A3",  X"BF",  X"2B",
  X"10",  X"C3",  X"10",  X"02",  X"3F",  X"0A",  X"0A",  X"32",
  X"12",  X"00",  X"12",  X"0A",  X"2A",  X"12",  X"0A",  X"C3",
  X"10",  X"10",  X"C3",  X"00",  X"E3",  X"10",  X"14",  X"04",
  X"A0",  X"80",  X"04",  X"C0",  X"04",  X"04",  X"A0",  X"BF",
  X"00",  X"C7",  X"E8",  X"E3",  X"C7",  X"E8",  X"00",  X"00",
  X"00",  X"00",  X"7A",  X"7C",  X"0C",  X"00",  X"00",  X"FF",
  X"00",  X"00",  X"00",  X"00",  X"7A",  X"04",  X"00",  X"98",
  X"00",  X"00",  X"00",  X"FF",  X"00",  X"41",  X"4E",  X"00",
  X"00",  X"00",  X"FF",  X"00",  X"41",  X"42",  X"00",  X"00",
  X"00",  X"FF",  X"00",  X"41",  X"46",  X"00",  X"00",  X"00",
  X"FF",  X"00",  X"41",  X"50",  X"00",  X"00",  X"00",  X"FF",
  X"00",  X"41",  X"57",  X"00",  X"00",  X"00",  X"FF",  X"00",
  X"41",  X"50",  X"00",  X"00",  X"00",  X"FF",  X"00",  X"41",
  X"4F",  X"00",  X"00",  X"00",  X"FF",  X"00",  X"41",  X"52",
  X"00",  X"00",  X"00",  X"FF",  X"00",  X"41",  X"50",  X"00",
  X"00",  X"00",  X"FF",  X"00",  X"41",  X"43",  X"00",  X"00",
  X"00",  X"FF",  X"00",  X"41",  X"42",  X"00",  X"00",  X"00",
  X"FF",  X"00",  X"00",  X"00",  X"00",  X"FF",  X"00",  X"41",
  X"4D",  X"00",  X"00",  X"00",  X"FF",  X"00",  X"41",  X"4E",
  X"00",  X"00",  X"00",  X"FF",  X"00",  X"41",  X"41",  X"00",
  X"00",  X"00",  X"FF",  X"00",  X"00",  X"00",  X"00",  X"FF",
  X"00",  X"00",  X"00",  X"00",  X"FF",  X"00",  X"41",  X"4C",
  X"00",  X"00",  X"00",  X"FF",  X"00",  X"00",  X"00",  X"00",
  X"FF",  X"00",  X"00",  X"00",  X"00",  X"FF",  X"00",  X"41",
  X"42",  X"00",  X"00",  X"00",  X"FF",  X"00",  X"41",  X"47",
  X"00",  X"00",  X"00",  X"FF",  X"00",  X"41",  X"09",  X"00",
  X"00",  X"FF",  X"00",  X"00",  X"00",  X"00",  X"FF",  X"00",
  X"41",  X"46",  X"00",  X"00",  X"00",  X"FF",  X"00",  X"00",
  X"00",  X"00",  X"FF",  X"00",  X"41",  X"4D",  X"00",  X"00",
  X"00",  X"FF",  X"00",  X"00",  X"00",  X"00",  X"FF",  X"00",
  X"41",  X"41",  X"00",  X"00",  X"00",  X"FF",  X"00",  X"41",
  X"49",  X"00",  X"00",  X"00",  X"FF",  X"00",  X"41",  X"4E",
  X"00",  X"00",  X"00",  X"FF",  X"00",  X"41",  X"51",  X"00",
  X"00",  X"00",  X"FF",  X"00",  X"41",  X"47",  X"00",  X"00",
  X"00",  X"FF",  X"00",  X"00",  X"00",  X"00",  X"FF",  X"00",
  X"00",  X"00",  X"00",  X"FF",  X"00",  X"41",  X"44",  X"00",
  X"00",  X"00",  X"FF",  X"00",  X"00",  X"00",  X"00",  X"FF",
  X"00",  X"41",  X"43",  X"00",  X"00",  X"00",  X"FF",  X"00",
  X"41",  X"44",  X"00",  X"00",  X"00",  X"FF",  X"00",  X"00",
  X"00",  X"00",  X"FF",  X"00",  X"41",  X"09",  X"00",  X"00",
  X"FF",  X"00",  X"41",  X"56",  X"00",  X"00",  X"00",  X"FF",
  X"00",  X"41",  X"4D",  X"00",  X"00",  X"00",  X"FF",  X"00",
  X"41",  X"46",  X"00",  X"00",  X"00",  X"FF",  X"00",  X"41",
  X"09",  X"00",  X"00",  X"FF",  X"00",  X"41",  X"09",  X"00",
  X"00",  X"FF",  X"00",  X"41",  X"43",  X"00",  X"00",  X"00",
  X"FF",  X"00",  X"41",  X"59",  X"00",  X"00",  X"00",  X"FF",
  X"00",  X"41",  X"09",  X"00",  X"00",  X"FF",  X"00",  X"41",
  X"09",  X"00",  X"00",  X"FF",  X"00",  X"00",  X"00",  X"00",
  X"FF",  X"00",  X"00",  X"00",  X"00",  X"FF",  X"00",  X"00",
  X"00",  X"00",  X"FF",  X"00",  X"41",  X"47",  X"00",  X"00",
  X"00",  X"FF",  X"00",  X"00",  X"00",  X"00",  X"FF",  X"00",
  X"41",  X"49",  X"00",  X"00",  X"00",  X"FF",  X"00",  X"41",
  X"5B",  X"00",  X"00",  X"00",  X"FF",  X"00",  X"41",  X"54",
  X"00",  X"00",  X"00",  X"FF",  X"00",  X"41",  X"56",  X"00",
  X"00",  X"00",  X"FF",  X"00",  X"41",  X"76",  X"00",  X"00",
  X"00",  X"FF",  X"00",  X"00",  X"00",  X"00",  X"FF",  X"00",
  X"00",  X"00",  X"00",  X"FF",  X"00",  X"00",  X"00",  X"00",
  X"FF",  X"00",  X"41",  X"57",  X"00",  X"00",  X"00",  X"FF",
  X"00",  X"45",  X"00",  X"00",  X"FF",  X"00",  X"41",  X"44",
  X"00",  X"00",  X"00",  X"FF",  X"00",  X"41",  X"41",  X"00",
  X"00",  X"00",  X"FF",  X"00",  X"00",  X"00",  X"00",  X"FF",
  X"00",  X"41",  X"4F",  X"00",  X"00",  X"00",  X"FF",  X"00",
  X"41",  X"43",  X"00",  X"00",  X"00",  X"FF",  X"00",  X"41",
  X"4A",  X"00",  X"00",  X"00",  X"FF",  X"00",  X"41",  X"4D",
  X"00",  X"00",  X"00",  X"FF",  X"00",  X"41",  X"4E",  X"00",
  X"00",  X"00",  X"FF",  X"00",  X"41",  X"41",  X"00",  X"00",
  X"00",  X"FF",  X"00",  X"41",  X"47",  X"00",  X"00",  X"00",
  X"FF",  X"00",  X"41",  X"47",  X"00",  X"00",  X"00",  X"FF",
  X"00",  X"41",  X"41",  X"00",  X"00",  X"00",  X"FF",  X"00",
  X"41",  X"43",  X"00",  X"00",  X"00",  X"FF",  X"00",  X"41",
  X"4F",  X"00",  X"00",  X"00",  X"FF",  X"00",  X"41",  X"44",
  X"00",  X"00",  X"00",  X"FF",  X"00",  X"41",  X"45",  X"00",
  X"00",  X"00",  X"FF",  X"00",  X"00",  X"00",  X"00",  X"FF",
  X"00",  X"00",  X"00",  X"00",  X"FF",  X"00",  X"00",  X"00",
  X"00",  X"FF",  X"00",  X"41",  X"44",  X"00",  X"00",  X"00",
  X"FF",  X"00",  X"41",  X"4A",  X"00",  X"00",  X"00",  X"FF",
  X"00",  X"41",  X"44",  X"00",  X"00",  X"00",  X"FF",  X"00",
  X"00",  X"00",  X"00",  X"FF",  X"00",  X"41",  X"5D",  X"00",
  X"00",  X"00",  X"FF",  X"00",  X"41",  X"44",  X"00",  X"00",
  X"00",  X"FF",  X"00",  X"41",  X"41",  X"00",  X"00",  X"00",
  X"FF",  X"00",  X"41",  X"42",  X"00",  X"00",  X"00",  X"FF",
  X"00",  X"41",  X"43",  X"00",  X"00",  X"00",  X"FF",  X"00",
  X"00",  X"00",  X"00",  X"FF",  X"00",  X"41",  X"43",  X"00",
  X"00",  X"00",  X"FF",  X"00",  X"41",  X"44",  X"00",  X"00",
  X"00",  X"FF",  X"00",  X"41",  X"44",  X"00",  X"00",  X"00",
  X"FF",  X"00",  X"00",  X"00",  X"00",  X"FF",  X"00",  X"00",
  X"00",  X"00",  X"FF",  X"00",  X"00",  X"00",  X"00",  X"FF",
  X"00",  X"41",  X"09",  X"00",  X"00",  X"FF",  X"00",  X"41",
  X"44",  X"00",  X"00",  X"00",  X"FF",  X"00",  X"00",  X"00",
  X"00",  X"FF",  X"00",  X"41",  X"45",  X"00",  X"00",  X"00",
  X"FF",  X"00",  X"00",  X"00",  X"00",  X"FF",  X"00",  X"00",
  X"00",  X"00",  X"FF",  X"00",  X"41",  X"52",  X"00",  X"00",
  X"00",  X"FF",  X"00",  X"00",  X"00",  X"00",  X"FF",  X"00",
  X"41",  X"58",  X"00",  X"00",  X"00",  X"FF",  X"00",  X"00",
  X"00",  X"00",  X"FF",  X"00",  X"41",  X"47",  X"00",  X"00",
  X"00",  X"FF",  X"00",  X"41",  X"45",  X"00",  X"00",  X"00",
  X"FF",  X"00",  X"41",  X"45",  X"00",  X"00",  X"00",  X"FF",
  X"00",  X"41",  X"45",  X"00",  X"00",  X"00",  X"FF",  X"00",
  X"41",  X"45",  X"00",  X"00",  X"00",  X"FF",  X"00",  X"41",
  X"45",  X"00",  X"00",  X"00",  X"FF",  X"00",  X"41",  X"45",
  X"00",  X"00",  X"00",  X"FF",  X"00",  X"41",  X"47",  X"00",
  X"00",  X"00",  X"FF",  X"00",  X"41",  X"47",  X"00",  X"00",
  X"00",  X"FF",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"FF",  X"00",  X"00",  X"00",  X"FF",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"73",  X"69",  X"52",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"09",  X"EB",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"31",  X"35",
  X"39",  X"44",  X"00",  X"00",  X"6E",  X"00",  X"31",  X"35",
  X"39",  X"64",  X"00",  X"00",  X"61",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"6E",  X"29",  X"00",  X"00",  X"30",  X"30",
  X"30",  X"30",  X"20",  X"20",  X"20",  X"20",  X"2D",  X"2D",
  X"2D",  X"53",  X"2D",  X"4A",  X"2D",  X"00",  X"6E",  X"69",
  X"00",  X"00",  X"F0",  X"00",  X"F8",  X"00",  X"D2",  X"6F",
  X"C6",  X"60",  X"D3",  X"9F",  X"F0",  X"00",  X"24",  X"00",
  X"1C",  X"00",  X"14",  X"00",  X"E0",  X"00",  X"53",  X"38",
  X"31",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"7F",  X"7F",  X"00",  X"00",
  X"F0",  X"00",  X"24",  X"00",  X"59",  X"00",  X"8F",  X"00",
  X"C3",  X"00",  X"F8",  X"00",  X"2E",  X"00",  X"63",  X"00",
  X"97",  X"00",  X"CD",  X"00",  X"02",  X"00",  X"37",  X"00",
  X"6D",  X"00",  X"A2",  X"40",  X"D6",  X"90",  X"0C",  X"34",
  X"41",  X"E0",  X"76",  X"D8",  X"AB",  X"4E",  X"E1",  X"91",
  X"15",  X"B5",  X"4B",  X"E2",  X"80",  X"4D",  X"B5",  X"E1",
  X"EA",  X"D9",  X"41",  X"E0",  X"93",  X"05",  X"38",  X"3F",
  X"82",  X"30",  X"15",  X"73",  X"9C",  X"D8",  X"49",  X"A8",
  X"A5",  X"F4",  X"5B",  X"8C",  X"C8",  X"AC",  X"00",  X"00",
  X"00",  X"00",  X"E3",  X"FF",  X"00",  X"FF",  X"00",  X"C7",
  X"E8",  X"E3",  X"FF",  X"00",  X"C7",  X"E8",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"0E",  X"34",  X"EC",  X"0B",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"02",  X"FF",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"FF",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  others => X"00" );


constant ram03 : ram_type := (
  X"88",  X"09",  X"81",  X"01",  X"A1",  X"A7",  X"10",  X"AC",
  X"91",  X"01",  X"01",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"A1",  X"29",  X"81",  X"01",  X"A1",  X"29",  X"81",  X"01",
  X"A1",  X"29",  X"81",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"91",  X"01",  X"01",  X"01",  X"A1",  X"A7",  X"10",  X"AC",
  X"91",  X"01",  X"01",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"91",  X"01",  X"01",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"91",  X"01",  X"01",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"91",  X"01",  X"01",  X"01",  X"AE",  X"A1",  X"10",  X"A7",
  X"AE",  X"A1",  X"10",  X"A7",  X"AE",  X"A1",  X"10",  X"A7",
  X"AE",  X"A1",  X"10",  X"A7",  X"AE",  X"A1",  X"10",  X"A7",
  X"AE",  X"A1",  X"10",  X"A7",  X"AE",  X"A1",  X"10",  X"A7",
  X"AE",  X"A1",  X"10",  X"A7",  X"AE",  X"A1",  X"10",  X"A7",
  X"AE",  X"A1",  X"10",  X"A7",  X"AE",  X"A1",  X"10",  X"A7",
  X"AE",  X"A1",  X"10",  X"A7",  X"AE",  X"A1",  X"10",  X"A7",
  X"AE",  X"A1",  X"10",  X"A7",  X"AE",  X"A1",  X"10",  X"A7",
  X"91",  X"01",  X"01",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"91",  X"01",  X"01",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"91",  X"01",  X"01",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"91",  X"01",  X"01",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"91",  X"01",  X"01",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"91",  X"01",  X"01",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"91",  X"01",  X"01",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"91",  X"01",  X"01",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"91",  X"01",  X"01",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"91",  X"01",  X"01",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"91",  X"01",  X"01",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"91",  X"01",  X"01",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"91",  X"01",  X"01",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"91",  X"01",  X"01",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"91",  X"01",  X"01",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"91",  X"01",  X"01",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"91",  X"01",  X"01",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"91",  X"01",  X"01",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"91",  X"01",  X"01",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"91",  X"01",  X"01",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"91",  X"01",  X"01",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"91",  X"01",  X"01",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"91",  X"01",  X"01",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"91",  X"01",  X"01",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"91",  X"01",  X"01",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"91",  X"01",  X"01",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"91",  X"01",  X"01",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"91",  X"01",  X"01",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"91",  X"01",  X"01",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"91",  X"01",  X"01",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"91",  X"01",  X"01",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"91",  X"01",  X"01",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"91",  X"01",  X"01",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"91",  X"01",  X"01",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"91",  X"01",  X"01",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"91",  X"01",  X"01",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"91",  X"01",  X"01",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"91",  X"01",  X"01",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"91",  X"01",  X"01",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"91",  X"01",  X"01",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"91",  X"01",  X"01",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"91",  X"01",  X"01",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"91",  X"01",  X"01",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"91",  X"01",  X"01",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"91",  X"01",  X"01",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"91",  X"01",  X"01",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"91",  X"01",  X"01",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"91",  X"01",  X"01",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"91",  X"01",  X"01",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"A1",  X"29",  X"81",  X"01",  X"A1",  X"10",  X"A7",  X"01",
  X"91",  X"01",  X"01",  X"01",  X"A1",  X"29",  X"81",  X"01",
  X"91",  X"01",  X"01",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"91",  X"01",  X"01",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"91",  X"01",  X"01",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"91",  X"01",  X"01",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"91",  X"01",  X"01",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"91",  X"01",  X"01",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"91",  X"01",  X"01",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"91",  X"01",  X"01",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"91",  X"01",  X"01",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"91",  X"01",  X"01",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"91",  X"01",  X"01",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"91",  X"01",  X"01",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"91",  X"01",  X"01",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"91",  X"01",  X"01",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"91",  X"01",  X"01",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"91",  X"01",  X"01",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"91",  X"01",  X"01",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"91",  X"01",  X"01",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"91",  X"01",  X"01",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"91",  X"01",  X"01",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"91",  X"01",  X"01",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"91",  X"01",  X"01",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"91",  X"01",  X"01",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"91",  X"01",  X"01",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"91",  X"01",  X"01",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"91",  X"01",  X"01",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"91",  X"01",  X"01",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"91",  X"01",  X"01",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"91",  X"01",  X"01",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"91",  X"01",  X"01",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"91",  X"01",  X"01",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"91",  X"01",  X"01",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"91",  X"01",  X"01",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"91",  X"01",  X"01",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"91",  X"01",  X"01",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"91",  X"01",  X"01",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"91",  X"01",  X"01",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"91",  X"01",  X"01",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"91",  X"01",  X"01",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"91",  X"01",  X"01",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"91",  X"01",  X"01",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"91",  X"01",  X"01",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"91",  X"01",  X"01",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"91",  X"01",  X"01",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"91",  X"01",  X"01",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"91",  X"01",  X"01",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"91",  X"01",  X"01",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"91",  X"01",  X"01",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"91",  X"01",  X"01",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"91",  X"01",  X"01",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"91",  X"01",  X"01",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"91",  X"01",  X"01",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"91",  X"01",  X"01",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"91",  X"01",  X"01",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"91",  X"01",  X"01",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"91",  X"01",  X"01",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"91",  X"01",  X"01",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"91",  X"01",  X"01",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"91",  X"01",  X"01",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"91",  X"01",  X"01",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"91",  X"01",  X"01",  X"01",  X"91",  X"01",  X"01",  X"01",
  X"9D",  X"05",  X"84",  X"07",  X"86",  X"82",  X"86",  X"86",
  X"36",  X"C0",  X"11",  X"90",  X"C0",  X"40",  X"01",  X"40",
  X"01",  X"40",  X"01",  X"11",  X"90",  X"40",  X"01",  X"40",
  X"01",  X"40",  X"01",  X"40",  X"01",  X"81",  X"81",  X"9D",
  X"21",  X"C2",  X"80",  X"12",  X"23",  X"C2",  X"27",  X"25",
  X"A6",  X"A4",  X"A4",  X"A5",  X"A4",  X"80",  X"3A",  X"03",
  X"A2",  X"82",  X"85",  X"C2",  X"C2",  X"9F",  X"01",  X"C2",
  X"80",  X"0A",  X"82",  X"03",  X"82",  X"80",  X"02",  X"82",
  X"11",  X"6F",  X"90",  X"82",  X"C2",  X"81",  X"81",  X"9D",
  X"81",  X"81",  X"9D",  X"03",  X"82",  X"80",  X"22",  X"11",
  X"11",  X"13",  X"90",  X"6F",  X"92",  X"11",  X"C2",  X"80",
  X"02",  X"90",  X"03",  X"82",  X"80",  X"02",  X"01",  X"9F",
  X"01",  X"81",  X"81",  X"9D",  X"81",  X"81",  X"81",  X"01",
  X"9D",  X"F2",  X"F4",  X"F6",  X"F8",  X"FA",  X"F0",  X"C0",
  X"82",  X"C2",  X"C2",  X"05",  X"90",  X"D2",  X"94",  X"40",
  X"01",  X"82",  X"C2",  X"03",  X"90",  X"03",  X"92",  X"D4",
  X"40",  X"01",  X"C2",  X"B0",  X"81",  X"81",  X"01",  X"9D",
  X"03",  X"90",  X"40",  X"01",  X"81",  X"81",  X"01",  X"9D",
  X"F0",  X"C2",  X"C2",  X"80",  X"12",  X"01",  X"C2",  X"C2",
  X"C4",  X"C4",  X"C6",  X"05",  X"84",  X"84",  X"C4",  X"10",
  X"01",  X"C2",  X"C2",  X"C4",  X"C6",  X"C4",  X"C4",  X"84",
  X"84",  X"C4",  X"85",  X"85",  X"C4",  X"C2",  X"C2",  X"84",
  X"C2",  X"C4",  X"C2",  X"C2",  X"82",  X"80",  X"82",  X"82",
  X"80",  X"02",  X"01",  X"C2",  X"C2",  X"C4",  X"C4",  X"C6",
  X"05",  X"84",  X"84",  X"C4",  X"10",  X"01",  X"C2",  X"C2",
  X"C2",  X"82",  X"82",  X"80",  X"82",  X"82",  X"80",  X"12",
  X"01",  X"81",  X"81",  X"01",  X"9D",  X"F0",  X"F2",  X"F4",
  X"C2",  X"C2",  X"C2",  X"C4",  X"C2",  X"84",  X"C2",  X"C4",
  X"C2",  X"C2",  X"80",  X"04",  X"01",  X"C2",  X"84",  X"C4",
  X"C0",  X"10",  X"01",  X"C2",  X"C4",  X"C2",  X"C2",  X"82",
  X"C6",  X"C8",  X"86",  X"C6",  X"C6",  X"C2",  X"C2",  X"C2",
  X"C2",  X"84",  X"C2",  X"C4",  X"C2",  X"C4",  X"C2",  X"82",
  X"80",  X"82",  X"82",  X"80",  X"02",  X"01",  X"C2",  X"84",
  X"C2",  X"C4",  X"C2",  X"82",  X"C2",  X"82",  X"C6",  X"C4",
  X"80",  X"06",  X"01",  X"82",  X"82",  X"80",  X"12",  X"01",
  X"C2",  X"C2",  X"80",  X"02",  X"01",  X"C2",  X"C2",  X"C4",
  X"C4",  X"C4",  X"86",  X"05",  X"84",  X"C4",  X"D0",  X"7F",
  X"01",  X"81",  X"81",  X"01",  X"9D",  X"F0",  X"C2",  X"05",
  X"84",  X"C4",  X"C2",  X"C2",  X"84",  X"C4",  X"C2",  X"84",
  X"C2",  X"C4",  X"C2",  X"C0",  X"C2",  X"C2",  X"05",  X"84",
  X"C4",  X"81",  X"81",  X"01",  X"9D",  X"F0",  X"C2",  X"05",
  X"84",  X"C4",  X"C2",  X"C2",  X"84",  X"C4",  X"C2",  X"C2",
  X"84",  X"C4",  X"C0",  X"10",  X"01",  X"C2",  X"C4",  X"C2",
  X"83",  X"82",  X"C0",  X"C2",  X"82",  X"C2",  X"82",  X"C4",
  X"80",  X"04",  X"01",  X"82",  X"82",  X"80",  X"12",  X"01",
  X"C2",  X"C2",  X"05",  X"84",  X"C4",  X"C2",  X"C2",  X"84",
  X"C4",  X"81",  X"81",  X"01",  X"9D",  X"03",  X"82",  X"C2",
  X"84",  X"03",  X"82",  X"C4",  X"03",  X"82",  X"C2",  X"05",
  X"90",  X"05",  X"92",  X"94",  X"7F",  X"01",  X"81",  X"81",
  X"01",  X"9D",  X"F0",  X"C2",  X"05",  X"84",  X"C4",  X"C2",
  X"C2",  X"C0",  X"C2",  X"C2",  X"C0",  X"C2",  X"C2",  X"84",
  X"C4",  X"03",  X"90",  X"92",  X"40",  X"01",  X"03",  X"90",
  X"92",  X"40",  X"01",  X"C2",  X"C2",  X"C4",  X"C4",  X"C4",
  X"84",  X"C4",  X"C2",  X"C2",  X"C4",  X"C4",  X"C4",  X"84",
  X"C4",  X"81",  X"81",  X"01",  X"9D",  X"F0",  X"F2",  X"C2",
  X"C2",  X"C4",  X"C4",  X"C6",  X"88",  X"C4",  X"85",  X"84",
  X"84",  X"C4",  X"81",  X"81",  X"01",  X"9D",  X"F0",  X"03",
  X"90",  X"7F",  X"01",  X"C2",  X"82",  X"90",  X"7F",  X"01",
  X"C2",  X"90",  X"7F",  X"01",  X"81",  X"81",  X"01",  X"9D",
  X"03",  X"90",  X"7F",  X"01",  X"03",  X"82",  X"C4",  X"C4",
  X"82",  X"C2",  X"10",  X"01",  X"92",  X"94",  X"90",  X"96",
  X"82",  X"40",  X"9E",  X"01",  X"9D",  X"82",  X"C2",  X"03",
  X"82",  X"C2",  X"C2",  X"82",  X"F2",  X"C2",  X"90",  X"F2",
  X"94",  X"96",  X"40",  X"92",  X"C2",  X"C0",  X"81",  X"91",
  X"9D",  X"03",  X"D0",  X"82",  X"C2",  X"03",  X"82",  X"C2",
  X"C2",  X"82",  X"F0",  X"F0",  X"C2",  X"94",  X"96",  X"40",
  X"92",  X"C2",  X"C0",  X"81",  X"91",  X"9D",  X"21",  X"40",
  X"90",  X"03",  X"E2",  X"D0",  X"80",  X"22",  X"90",  X"C2",
  X"80",  X"14",  X"01",  X"80",  X"02",  X"84",  X"C4",  X"82",
  X"86",  X"89",  X"87",  X"C2",  X"F4",  X"F6",  X"86",  X"87",
  X"82",  X"C2",  X"80",  X"02",  X"82",  X"84",  X"85",  X"82",
  X"C2",  X"F2",  X"B0",  X"40",  X"90",  X"81",  X"81",  X"40",
  X"90",  X"80",  X"22",  X"90",  X"C2",  X"C2",  X"D0",  X"C0",
  X"C0",  X"C0",  X"10",  X"82",  X"C2",  X"86",  X"82",  X"84",
  X"85",  X"C6",  X"82",  X"F2",  X"C2",  X"B0",  X"40",  X"90",
  X"81",  X"81",  X"10",  X"D0",  X"40",  X"B0",  X"81",  X"81",
  X"92",  X"03",  X"D0",  X"82",  X"40",  X"9E",  X"01",  X"92",
  X"03",  X"D0",  X"82",  X"40",  X"9E",  X"01",  X"9D",  X"84",
  X"82",  X"80",  X"08",  X"A0",  X"A0",  X"85",  X"80",  X"0A",
  X"80",  X"12",  X"01",  X"40",  X"90",  X"80",  X"18",  X"83",
  X"23",  X"A2",  X"82",  X"E4",  X"80",  X"02",  X"99",  X"C6",
  X"C4",  X"C2",  X"86",  X"86",  X"C8",  X"88",  X"C2",  X"C8",
  X"C4",  X"90",  X"40",  X"B0",  X"81",  X"81",  X"E6",  X"E8",
  X"A8",  X"82",  X"80",  X"14",  X"80",  X"03",  X"2F",  X"EA",
  X"C2",  X"AA",  X"80",  X"02",  X"AA",  X"AA",  X"AA",  X"90",
  X"40",  X"92",  X"80",  X"02",  X"A4",  X"84",  X"80",  X"08",
  X"2D",  X"80",  X"02",  X"C2",  X"C2",  X"C4",  X"84",  X"82",
  X"80",  X"14",  X"80",  X"40",  X"90",  X"81",  X"91",  X"99",
  X"80",  X"02",  X"87",  X"80",  X"08",  X"99",  X"98",  X"80",
  X"08",  X"87",  X"80",  X"18",  X"80",  X"99",  X"98",  X"87",
  X"23",  X"A2",  X"86",  X"E4",  X"80",  X"32",  X"C4",  X"10",
  X"98",  X"36",  X"C6",  X"E4",  X"80",  X"22",  X"98",  X"C4",
  X"84",  X"82",  X"80",  X"04",  X"80",  X"98",  X"98",  X"07",
  X"86",  X"E4",  X"80",  X"22",  X"C2",  X"C4",  X"84",  X"82",
  X"80",  X"14",  X"80",  X"C6",  X"16",  X"C6",  X"80",  X"28",
  X"85",  X"83",  X"80",  X"18",  X"88",  X"89",  X"88",  X"9B",
  X"9A",  X"C2",  X"80",  X"32",  X"C8",  X"10",  X"DA",  X"80",
  X"22",  X"C4",  X"C8",  X"88",  X"80",  X"2A",  X"C2",  X"C4",
  X"C4",  X"C2",  X"E4",  X"E4",  X"C2",  X"85",  X"88",  X"89",
  X"80",  X"2A",  X"E6",  X"80",  X"22",  X"98",  X"95",  X"96",
  X"94",  X"9A",  X"E4",  X"80",  X"32",  X"C4",  X"10",  X"96",
  X"36",  X"C6",  X"E4",  X"80",  X"22",  X"96",  X"C4",  X"84",
  X"82",  X"80",  X"04",  X"80",  X"DA",  X"C8",  X"84",  X"A0",
  X"C8",  X"DA",  X"C4",  X"C4",  X"E0",  X"C2",  X"C6",  X"10",
  X"C6",  X"C2",  X"84",  X"C8",  X"88",  X"C2",  X"C8",  X"C6",
  X"90",  X"40",  X"B0",  X"81",  X"81",  X"84",  X"C2",  X"82",
  X"C2",  X"90",  X"40",  X"B0",  X"81",  X"81",  X"98",  X"10",
  X"87",  X"89",  X"88",  X"DA",  X"D6",  X"C8",  X"DA",  X"85",
  X"82",  X"E4",  X"83",  X"E4",  X"82",  X"10",  X"C2",  X"89",
  X"80",  X"02",  X"98",  X"10",  X"95",  X"38",  X"03",  X"E4",
  X"84",  X"A0",  X"82",  X"E0",  X"C2",  X"90",  X"C4",  X"40",
  X"B0",  X"81",  X"81",  X"84",  X"10",  X"A0",  X"80",  X"12",
  X"9A",  X"80",  X"02",  X"82",  X"D4",  X"80",  X"22",  X"98",
  X"C2",  X"89",  X"80",  X"18",  X"80",  X"22",  X"E6",  X"80",
  X"22",  X"89",  X"10",  X"98",  X"82",  X"E4",  X"80",  X"02",
  X"98",  X"10",  X"C6",  X"C2",  X"82",  X"80",  X"02",  X"C2",
  X"C6",  X"80",  X"22",  X"03",  X"82",  X"84",  X"C4",  X"84",
  X"02",  X"03",  X"82",  X"82",  X"A4",  X"82",  X"AA",  X"90",
  X"AA",  X"AA",  X"40",  X"92",  X"80",  X"02",  X"84",  X"84",
  X"84",  X"84",  X"C2",  X"82",  X"C2",  X"C4",  X"80",  X"02",
  X"E4",  X"80",  X"08",  X"84",  X"84",  X"86",  X"C8",  X"88",
  X"88",  X"C8",  X"88",  X"C8",  X"80",  X"18",  X"C8",  X"05",
  X"C6",  X"80",  X"38",  X"C2",  X"05",  X"C6",  X"80",  X"38",
  X"C2",  X"10",  X"C2",  X"28",  X"E4",  X"30",  X"18",  X"80",
  X"99",  X"98",  X"10",  X"87",  X"80",  X"08",  X"9B",  X"80",
  X"18",  X"80",  X"89",  X"88",  X"10",  X"9B",  X"89",  X"84",
  X"85",  X"84",  X"C4",  X"10",  X"84",  X"86",  X"18",  X"98",
  X"99",  X"98",  X"10",  X"87",  X"82",  X"10",  X"C2",  X"18",
  X"80",  X"89",  X"88",  X"10",  X"9B",  X"80",  X"12",  X"C6",
  X"C4",  X"86",  X"86",  X"10",  X"C6",  X"10",  X"E4",  X"92",
  X"40",  X"90",  X"03",  X"10",  X"C2",  X"10",  X"AA",  X"9A",
  X"18",  X"88",  X"89",  X"88",  X"10",  X"9B",  X"C2",  X"82",
  X"10",  X"C2",  X"10",  X"96",  X"11",  X"90",  X"82",  X"40",
  X"9E",  X"01",  X"11",  X"90",  X"82",  X"40",  X"9E",  X"01",
  X"9D",  X"21",  X"90",  X"40",  X"C0",  X"80",  X"02",  X"C2",
  X"81",  X"91",  X"80",  X"02",  X"01",  X"C2",  X"81",  X"91",
  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",
  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",
  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",
  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",
  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",
  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",
  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",
  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",
  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",
  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",
  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",
  X"40",  X"9D",  X"C2",  X"80",  X"12",  X"90",  X"C0",  X"81",
  X"91",  X"40",  X"92",  X"C0",  X"C0",  X"81",  X"91",  X"9D",
  X"40",  X"01",  X"D0",  X"C2",  X"F0",  X"80",  X"02",  X"D0",
  X"03",  X"D0",  X"80",  X"22",  X"C2",  X"C2",  X"80",  X"02",
  X"01",  X"C2",  X"80",  X"02",  X"86",  X"C4",  X"80",  X"02",
  X"84",  X"80",  X"22",  X"C4",  X"A6",  X"C0",  X"C0",  X"E6",
  X"C0",  X"C0",  X"C0",  X"C0",  X"25",  X"23",  X"A4",  X"A2",
  X"B0",  X"A0",  X"C4",  X"80",  X"02",  X"C2",  X"80",  X"02",
  X"83",  X"A8",  X"A8",  X"C2",  X"80",  X"02",  X"80",  X"32",
  X"A8",  X"AA",  X"22",  X"B4",  X"EA",  X"F4",  X"A0",  X"C2",
  X"C4",  X"82",  X"84",  X"C2",  X"80",  X"14",  X"C4",  X"C2",
  X"B4",  X"B0",  X"83",  X"80",  X"02",  X"B4",  X"C0",  X"AC",
  X"EA",  X"AB",  X"B8",  X"A8",  X"86",  X"88",  X"AB",  X"B4",
  X"82",  X"80",  X"28",  X"83",  X"80",  X"02",  X"84",  X"EA",
  X"C0",  X"C4",  X"C0",  X"BA",  X"AE",  X"AC",  X"80",  X"02",
  X"86",  X"C4",  X"84",  X"C4",  X"02",  X"C6",  X"C2",  X"80",
  X"02",  X"80",  X"82",  X"C2",  X"82",  X"C2",  X"C4",  X"C2",
  X"82",  X"84",  X"C2",  X"C4",  X"80",  X"14",  X"A0",  X"C2",
  X"80",  X"02",  X"C4",  X"C4",  X"82",  X"80",  X"04",  X"80",
  X"04",  X"E2",  X"86",  X"84",  X"A0",  X"10",  X"82",  X"A0",
  X"80",  X"24",  X"84",  X"C4",  X"E2",  X"82",  X"C6",  X"C8",
  X"86",  X"88",  X"C6",  X"80",  X"04",  X"C8",  X"C4",  X"90",
  X"7F",  X"92",  X"80",  X"12",  X"C4",  X"A0",  X"80",  X"14",
  X"82",  X"84",  X"82",  X"A0",  X"C2",  X"C6",  X"C6",  X"C4",
  X"82",  X"C2",  X"C2",  X"82",  X"C2",  X"80",  X"04",  X"A0",
  X"90",  X"7F",  X"92",  X"80",  X"12",  X"A0",  X"80",  X"12",
  X"80",  X"FA",  X"EE",  X"A0",  X"C2",  X"BA",  X"FA",  X"C2",
  X"82",  X"80",  X"14",  X"C2",  X"80",  X"02",  X"E8",  X"C2",
  X"A8",  X"80",  X"04",  X"80",  X"04",  X"E4",  X"AA",  X"10",
  X"AE",  X"A8",  X"80",  X"24",  X"E8",  X"EA",  X"E4",  X"A0",
  X"C2",  X"C4",  X"82",  X"84",  X"C2",  X"80",  X"04",  X"C4",
  X"90",  X"7F",  X"92",  X"80",  X"12",  X"A8",  X"80",  X"14",
  X"A0",  X"E8",  X"C4",  X"C4",  X"C2",  X"A8",  X"C2",  X"82",
  X"E8",  X"80",  X"04",  X"C2",  X"90",  X"7F",  X"92",  X"80",
  X"12",  X"80",  X"E8",  X"C6",  X"80",  X"26",  X"B8",  X"80",
  X"12",  X"B0",  X"C0",  X"80",  X"02",  X"A0",  X"D0",  X"40",
  X"92",  X"10",  X"C4",  X"05",  X"84",  X"C2",  X"81",  X"01",
  X"10",  X"C2",  X"A8",  X"80",  X"32",  X"FA",  X"80",  X"22",
  X"FA",  X"FA",  X"80",  X"B6",  X"84",  X"82",  X"C0",  X"80",
  X"36",  X"A8",  X"86",  X"80",  X"12",  X"C6",  X"80",  X"02",
  X"80",  X"82",  X"80",  X"02",  X"80",  X"02",  X"AE",  X"82",
  X"AE",  X"82",  X"BB",  X"80",  X"12",  X"C2",  X"C4",  X"80",
  X"02",  X"BA",  X"80",  X"02",  X"82",  X"AE",  X"BA",  X"10",
  X"C2",  X"80",  X"B6",  X"84",  X"10",  X"82",  X"A8",  X"80",
  X"32",  X"FA",  X"80",  X"22",  X"FA",  X"FA",  X"80",  X"B6",
  X"84",  X"10",  X"82",  X"80",  X"B6",  X"84",  X"10",  X"82",
  X"A8",  X"80",  X"02",  X"80",  X"FA",  X"B6",  X"80",  X"06",
  X"80",  X"82",  X"10",  X"84",  X"12",  X"AE",  X"80",  X"12",
  X"82",  X"AE",  X"BA",  X"80",  X"16",  X"FA",  X"EC",  X"EC",
  X"AC",  X"C2",  X"80",  X"02",  X"80",  X"C2",  X"82",  X"C2",
  X"86",  X"12",  X"C6",  X"C4",  X"82",  X"80",  X"04",  X"80",
  X"04",  X"E4",  X"86",  X"84",  X"A0",  X"10",  X"82",  X"A0",
  X"80",  X"24",  X"84",  X"C4",  X"E4",  X"82",  X"C6",  X"C8",
  X"86",  X"88",  X"C6",  X"80",  X"04",  X"C8",  X"C4",  X"90",
  X"7F",  X"92",  X"80",  X"12",  X"C4",  X"A0",  X"80",  X"14",
  X"82",  X"84",  X"82",  X"A0",  X"C2",  X"C6",  X"C6",  X"C4",
  X"82",  X"C2",  X"C2",  X"82",  X"C2",  X"80",  X"04",  X"A0",
  X"90",  X"7F",  X"92",  X"80",  X"12",  X"C2",  X"80",  X"12",
  X"A0",  X"80",  X"02",  X"C2",  X"EA",  X"82",  X"C2",  X"82",
  X"C2",  X"82",  X"C2",  X"C4",  X"C2",  X"82",  X"84",  X"C2",
  X"C4",  X"80",  X"04",  X"A0",  X"90",  X"7F",  X"92",  X"80",
  X"12",  X"C2",  X"80",  X"12",  X"A0",  X"C4",  X"82",  X"80",
  X"04",  X"80",  X"04",  X"E2",  X"86",  X"84",  X"A0",  X"10",
  X"82",  X"A0",  X"80",  X"24",  X"84",  X"C4",  X"E2",  X"82",
  X"C6",  X"C8",  X"86",  X"88",  X"C6",  X"80",  X"04",  X"C8",
  X"C4",  X"90",  X"7F",  X"92",  X"80",  X"12",  X"C4",  X"A0",
  X"80",  X"14",  X"82",  X"84",  X"82",  X"A0",  X"C2",  X"C6",
  X"C6",  X"C4",  X"82",  X"C2",  X"C2",  X"82",  X"C2",  X"80",
  X"04",  X"A0",  X"90",  X"7F",  X"92",  X"80",  X"12",  X"A0",
  X"10",  X"C4",  X"04",  X"C2",  X"03",  X"D5",  X"82",  X"D1",
  X"81",  X"01",  X"03",  X"C2",  X"82",  X"C2",  X"03",  X"82",
  X"C4",  X"C2",  X"C2",  X"82",  X"84",  X"C2",  X"C4",  X"80",
  X"14",  X"A0",  X"C2",  X"C4",  X"80",  X"06",  X"82",  X"80",
  X"02",  X"80",  X"82",  X"C2",  X"C6",  X"C6",  X"C2",  X"C4",
  X"82",  X"84",  X"C2",  X"C4",  X"80",  X"14",  X"A0",  X"C2",
  X"AA",  X"80",  X"04",  X"80",  X"04",  X"E2",  X"AE",  X"10",
  X"BA",  X"AA",  X"80",  X"24",  X"EA",  X"EE",  X"E2",  X"A0",
  X"C2",  X"C4",  X"82",  X"84",  X"C2",  X"80",  X"04",  X"C4",
  X"90",  X"7F",  X"92",  X"80",  X"12",  X"A0",  X"10",  X"AA",
  X"90",  X"7F",  X"92",  X"80",  X"22",  X"C0",  X"80",  X"22",
  X"C2",  X"D0",  X"40",  X"92",  X"C2",  X"83",  X"83",  X"80",
  X"02",  X"01",  X"80",  X"12",  X"01",  X"81",  X"81",  X"81",
  X"91",  X"40",  X"90",  X"80",  X"32",  X"C2",  X"C6",  X"82",
  X"84",  X"80",  X"12",  X"A6",  X"C4",  X"80",  X"06",  X"C4",
  X"80",  X"02",  X"01",  X"86",  X"C2",  X"C2",  X"82",  X"C8",
  X"C2",  X"C2",  X"82",  X"C6",  X"C4",  X"C8",  X"A2",  X"C2",
  X"C2",  X"90",  X"40",  X"C0",  X"90",  X"40",  X"92",  X"92",
  X"A0",  X"40",  X"90",  X"40",  X"90",  X"D0",  X"A2",  X"94",
  X"92",  X"7F",  X"96",  X"B0",  X"06",  X"C2",  X"40",  X"90",
  X"80",  X"32",  X"B0",  X"C2",  X"80",  X"02",  X"01",  X"C2",
  X"82",  X"C2",  X"40",  X"90",  X"81",  X"81",  X"80",  X"04",
  X"80",  X"C2",  X"C2",  X"82",  X"C2",  X"82",  X"C2",  X"82",
  X"C2",  X"C4",  X"C2",  X"82",  X"84",  X"C2",  X"C4",  X"80",
  X"14",  X"A0",  X"05",  X"D5",  X"84",  X"D1",  X"81",  X"01",
  X"13",  X"C6",  X"C4",  X"82",  X"C2",  X"AE",  X"EE",  X"C4",
  X"82",  X"C2",  X"C2",  X"82",  X"C2",  X"80",  X"14",  X"A0",
  X"C4",  X"C4",  X"82",  X"C6",  X"C2",  X"C4",  X"C2",  X"82",
  X"84",  X"C4",  X"C2",  X"80",  X"04",  X"A0",  X"90",  X"7F",
  X"92",  X"80",  X"12",  X"A0",  X"10",  X"80",  X"90",  X"7F",
  X"92",  X"80",  X"12",  X"A0",  X"10",  X"C2",  X"40",  X"90",
  X"10",  X"03",  X"40",  X"01",  X"10",  X"C2",  X"40",  X"90",
  X"10",  X"C2",  X"80",  X"04",  X"C4",  X"80",  X"26",  X"C2",
  X"C4",  X"C6",  X"EE",  X"C2",  X"C4",  X"82",  X"84",  X"C2",
  X"C4",  X"80",  X"14",  X"A0",  X"EA",  X"C2",  X"AA",  X"80",
  X"04",  X"80",  X"04",  X"E2",  X"AE",  X"10",  X"BA",  X"AA",
  X"80",  X"24",  X"EA",  X"EE",  X"E2",  X"A0",  X"C2",  X"C4",
  X"82",  X"84",  X"C2",  X"80",  X"04",  X"C4",  X"90",  X"7F",
  X"92",  X"80",  X"12",  X"A0",  X"10",  X"AA",  X"AE",  X"C2",
  X"10",  X"BA",  X"AA",  X"80",  X"04",  X"80",  X"04",  X"E2",
  X"AE",  X"10",  X"BA",  X"AA",  X"80",  X"24",  X"EA",  X"EE",
  X"E2",  X"A0",  X"C2",  X"C4",  X"82",  X"84",  X"C2",  X"80",
  X"04",  X"C4",  X"90",  X"7F",  X"92",  X"80",  X"12",  X"A0",
  X"10",  X"AA",  X"22",  X"FA",  X"FA",  X"10",  X"B6",  X"40",
  X"90",  X"C6",  X"10",  X"C4",  X"F8",  X"80",  X"16",  X"B6",
  X"B8",  X"EA",  X"A8",  X"10",  X"AB",  X"80",  X"02",  X"80",
  X"32",  X"AC",  X"C2",  X"BA",  X"B6",  X"AE",  X"C2",  X"82",
  X"C0",  X"83",  X"C0",  X"82",  X"AC",  X"10",  X"C2",  X"80",
  X"12",  X"C2",  X"80",  X"02",  X"01",  X"B6",  X"10",  X"F0",
  X"EA",  X"A8",  X"10",  X"AB",  X"EA",  X"10",  X"AB",  X"C6",
  X"EA",  X"10",  X"AB",  X"EA",  X"A8",  X"10",  X"AB",  X"82",
  X"B8",  X"EA",  X"85",  X"B9",  X"B8",  X"B8",  X"82",  X"80",
  X"08",  X"B4",  X"10",  X"82",  X"FA",  X"80",  X"07",  X"B6",
  X"86",  X"84",  X"A8",  X"C6",  X"82",  X"10",  X"AA",  X"EA",
  X"A8",  X"10",  X"AB",  X"EA",  X"AB",  X"83",  X"80",  X"22",
  X"B4",  X"10",  X"A8",  X"03",  X"82",  X"80",  X"12",  X"C2",
  X"80",  X"22",  X"FA",  X"FA",  X"B6",  X"80",  X"84",  X"80",
  X"02",  X"82",  X"80",  X"22",  X"C0",  X"A8",  X"10",  X"84",
  X"EA",  X"80",  X"02",  X"B4",  X"82",  X"84",  X"80",  X"18",
  X"AC",  X"EA",  X"9B",  X"85",  X"84",  X"84",  X"82",  X"80",
  X"08",  X"B4",  X"AC",  X"26",  X"AC",  X"10",  X"82",  X"EA",
  X"A8",  X"10",  X"AB",  X"C0",  X"EE",  X"80",  X"02",  X"B6",
  X"80",  X"02",  X"80",  X"32",  X"EE",  X"80",  X"06",  X"90",
  X"92",  X"40",  X"94",  X"80",  X"22",  X"EC",  X"BA",  X"80",
  X"04",  X"82",  X"EC",  X"BA",  X"C0",  X"10",  X"AC",  X"07",
  X"86",  X"80",  X"02",  X"C6",  X"FA",  X"10",  X"B6",  X"C2",
  X"80",  X"32",  X"EA",  X"C8",  X"EA",  X"10",  X"AB",  X"EA",
  X"A8",  X"10",  X"AB",  X"80",  X"02",  X"80",  X"02",  X"80",
  X"02",  X"80",  X"80",  X"02",  X"92",  X"90",  X"40",  X"94",
  X"D1",  X"D1",  X"D1",  X"B6",  X"40",  X"D0",  X"80",  X"02",
  X"03",  X"D5",  X"82",  X"D1",  X"81",  X"01",  X"09",  X"82",
  X"82",  X"2F",  X"C2",  X"BA",  X"C0",  X"AE",  X"10",  X"AC",
  X"B6",  X"10",  X"F0",  X"C4",  X"82",  X"C2",  X"AE",  X"BB",
  X"80",  X"12",  X"C2",  X"C2",  X"10",  X"BA",  X"80",  X"08",
  X"84",  X"AE",  X"90",  X"92",  X"40",  X"AE",  X"82",  X"92",
  X"90",  X"40",  X"C2",  X"80",  X"18",  X"BA",  X"84",  X"82",
  X"C6",  X"AE",  X"C2",  X"10",  X"BA",  X"32",  X"C2",  X"82",
  X"C2",  X"EE",  X"A0",  X"C2",  X"C4",  X"82",  X"84",  X"C2",
  X"80",  X"04",  X"C4",  X"90",  X"7F",  X"92",  X"80",  X"12",
  X"A0",  X"10",  X"C4",  X"90",  X"7F",  X"92",  X"80",  X"12",
  X"A0",  X"10",  X"05",  X"EA",  X"C2",  X"C2",  X"C2",  X"AA",
  X"C2",  X"82",  X"EA",  X"C2",  X"80",  X"04",  X"A0",  X"10",
  X"90",  X"AC",  X"92",  X"94",  X"40",  X"90",  X"D4",  X"D0",
  X"96",  X"AE",  X"40",  X"92",  X"80",  X"02",  X"BA",  X"10",
  X"B6",  X"82",  X"BA",  X"C2",  X"80",  X"82",  X"10",  X"84",
  X"EA",  X"C4",  X"C4",  X"C2",  X"AA",  X"A0",  X"10",  X"EA",
  X"90",  X"40",  X"94",  X"D5",  X"D5",  X"B6",  X"10",  X"D5",
  X"EE",  X"92",  X"90",  X"40",  X"94",  X"80",  X"06",  X"BA",
  X"82",  X"F6",  X"B6",  X"AA",  X"A0",  X"BA",  X"10",  X"AC",
  X"A0",  X"C2",  X"D4",  X"80",  X"02",  X"D0",  X"92",  X"40",
  X"96",  X"80",  X"22",  X"C4",  X"82",  X"80",  X"14",  X"80",
  X"12",  X"AC",  X"A0",  X"AA",  X"F6",  X"80",  X"12",  X"AC",
  X"C0",  X"10",  X"C0",  X"EE",  X"A0",  X"C4",  X"82",  X"C2",
  X"C2",  X"82",  X"80",  X"14",  X"C2",  X"82",  X"EA",  X"C2",
  X"03",  X"82",  X"C4",  X"C2",  X"C2",  X"82",  X"84",  X"C2",
  X"C4",  X"80",  X"14",  X"A0",  X"C2",  X"C6",  X"84",  X"C4",
  X"AA",  X"EA",  X"C4",  X"84",  X"C2",  X"10",  X"82",  X"EA",
  X"C4",  X"C4",  X"C2",  X"AA",  X"C2",  X"82",  X"EA",  X"C2",
  X"80",  X"04",  X"A0",  X"90",  X"7F",  X"92",  X"80",  X"12",
  X"A0",  X"80",  X"02",  X"80",  X"82",  X"C2",  X"03",  X"82",
  X"C4",  X"C2",  X"C2",  X"82",  X"10",  X"84",  X"80",  X"22",
  X"AC",  X"10",  X"80",  X"90",  X"7F",  X"92",  X"80",  X"12",
  X"A0",  X"10",  X"C2",  X"84",  X"2F",  X"C2",  X"C4",  X"BA",
  X"AE",  X"C0",  X"10",  X"AC",  X"82",  X"C2",  X"03",  X"82",
  X"C4",  X"C2",  X"C2",  X"82",  X"84",  X"C2",  X"C4",  X"80",
  X"14",  X"A0",  X"C2",  X"80",  X"02",  X"C6",  X"82",  X"C2",
  X"C2",  X"C2",  X"C4",  X"C6",  X"84",  X"86",  X"C4",  X"C6",
  X"80",  X"14",  X"82",  X"EA",  X"AA",  X"80",  X"04",  X"80",
  X"04",  X"E2",  X"BA",  X"10",  X"A0",  X"AA",  X"80",  X"24",
  X"EA",  X"FA",  X"E2",  X"82",  X"C4",  X"C6",  X"84",  X"86",
  X"C4",  X"80",  X"04",  X"C6",  X"90",  X"7F",  X"92",  X"80",
  X"12",  X"82",  X"10",  X"AA",  X"80",  X"02",  X"80",  X"10",
  X"82",  X"90",  X"7F",  X"92",  X"80",  X"12",  X"A0",  X"10",
  X"EA",  X"90",  X"7F",  X"92",  X"80",  X"12",  X"A0",  X"10",
  X"C2",  X"90",  X"7F",  X"92",  X"80",  X"12",  X"A0",  X"10",
  X"82",  X"90",  X"7F",  X"92",  X"80",  X"12",  X"A0",  X"10",
  X"C2",  X"C0",  X"40",  X"AC",  X"82",  X"BA",  X"83",  X"82",
  X"10",  X"C2",  X"C2",  X"80",  X"12",  X"90",  X"C0",  X"10",
  X"C2",  X"7F",  X"92",  X"80",  X"32",  X"C2",  X"C0",  X"10",
  X"C2",  X"10",  X"AC",  X"EA",  X"A8",  X"10",  X"AB",  X"40",
  X"D0",  X"80",  X"12",  X"86",  X"A8",  X"80",  X"BA",  X"02",
  X"96",  X"80",  X"02",  X"80",  X"02",  X"96",  X"D1",  X"D1",
  X"C0",  X"C2",  X"80",  X"06",  X"95",  X"82",  X"D0",  X"C2",
  X"D2",  X"82",  X"D4",  X"C2",  X"98",  X"40",  X"9A",  X"80",
  X"02",  X"AE",  X"80",  X"02",  X"80",  X"03",  X"80",  X"84",
  X"02",  X"82",  X"D1",  X"D5",  X"81",  X"01",  X"03",  X"C8",
  X"C4",  X"82",  X"84",  X"80",  X"82",  X"80",  X"02",  X"C4",
  X"80",  X"02",  X"80",  X"FA",  X"80",  X"06",  X"80",  X"80",
  X"16",  X"C6",  X"80",  X"AA",  X"02",  X"82",  X"82",  X"AA",
  X"BA",  X"C2",  X"80",  X"06",  X"FA",  X"82",  X"C2",  X"80",
  X"14",  X"82",  X"BA",  X"82",  X"C2",  X"FA",  X"84",  X"C2",
  X"80",  X"82",  X"82",  X"C4",  X"C2",  X"04",  X"BA",  X"BA",
  X"C4",  X"80",  X"02",  X"82",  X"82",  X"C0",  X"C2",  X"AC",
  X"82",  X"83",  X"82",  X"82",  X"10",  X"C2",  X"80",  X"02",
  X"C4",  X"10",  X"BA",  X"90",  X"7F",  X"92",  X"80",  X"12",
  X"A0",  X"10",  X"C2",  X"C0",  X"83",  X"AC",  X"82",  X"10",
  X"C2",  X"EA",  X"C4",  X"C4",  X"C4",  X"AA",  X"C4",  X"84",
  X"EA",  X"C4",  X"80",  X"04",  X"82",  X"90",  X"7F",  X"92",
  X"80",  X"12",  X"82",  X"C6",  X"C6",  X"EE",  X"A0",  X"C4",
  X"C2",  X"82",  X"84",  X"C2",  X"80",  X"04",  X"C4",  X"10",
  X"90",  X"82",  X"2F",  X"C2",  X"BA",  X"AE",  X"C0",  X"10",
  X"AC",  X"2F",  X"C6",  X"BA",  X"C0",  X"AE",  X"10",  X"AC",
  X"D0",  X"7F",  X"92",  X"AC",  X"02",  X"94",  X"92",  X"40",
  X"90",  X"D0",  X"92",  X"98",  X"94",  X"40",  X"96",  X"80",
  X"12",  X"82",  X"C0",  X"AE",  X"83",  X"C0",  X"82",  X"10",
  X"C2",  X"80",  X"12",  X"90",  X"40",  X"B0",  X"81",  X"81",
  X"BA",  X"A0",  X"AA",  X"10",  X"F6",  X"04",  X"80",  X"02",
  X"FA",  X"C6",  X"80",  X"14",  X"80",  X"80",  X"02",  X"AA",
  X"10",  X"BA",  X"80",  X"12",  X"03",  X"10",  X"C4",  X"80",
  X"82",  X"08",  X"86",  X"C6",  X"82",  X"80",  X"18",  X"C2",
  X"10",  X"82",  X"D0",  X"92",  X"94",  X"96",  X"40",  X"98",
  X"80",  X"02",  X"BA",  X"10",  X"EE",  X"90",  X"7F",  X"92",
  X"80",  X"12",  X"82",  X"10",  X"EA",  X"C4",  X"84",  X"82",
  X"10",  X"C4",  X"BA",  X"10",  X"96",  X"AC",  X"C2",  X"90",
  X"92",  X"40",  X"AC",  X"84",  X"92",  X"90",  X"40",  X"C4",
  X"C2",  X"80",  X"14",  X"BA",  X"88",  X"84",  X"86",  X"C8",
  X"80",  X"18",  X"84",  X"10",  X"C2",  X"C8",  X"86",  X"C8",
  X"80",  X"18",  X"84",  X"10",  X"C2",  X"FA",  X"10",  X"82",
  X"97",  X"95",  X"82",  X"D5",  X"10",  X"C2",  X"C2",  X"80",
  X"02",  X"03",  X"FA",  X"84",  X"10",  X"82",  X"82",  X"04",
  X"BA",  X"BA",  X"C2",  X"BA",  X"10",  X"AA",  X"07",  X"D5",
  X"86",  X"D1",  X"81",  X"01",  X"13",  X"82",  X"86",  X"BA",
  X"FA",  X"10",  X"84",  X"82",  X"BA",  X"10",  X"C2",  X"FA",
  X"10",  X"84",  X"EC",  X"80",  X"16",  X"B6",  X"EA",  X"AB",
  X"10",  X"AC",  X"80",  X"04",  X"80",  X"32",  X"BA",  X"80",
  X"02",  X"C4",  X"BA",  X"AA",  X"10",  X"BA",  X"12",  X"BA",
  X"80",  X"02",  X"BA",  X"BA",  X"10",  X"AA",  X"10",  X"84",
  X"C2",  X"82",  X"10",  X"C2",  X"03",  X"84",  X"D0",  X"82",
  X"96",  X"92",  X"94",  X"82",  X"7F",  X"9E",  X"01",  X"9D",
  X"80",  X"02",  X"A0",  X"92",  X"94",  X"90",  X"40",  X"96",
  X"80",  X"12",  X"B0",  X"C0",  X"82",  X"C2",  X"81",  X"81",
  X"90",  X"92",  X"94",  X"40",  X"96",  X"10",  X"80",  X"03",
  X"84",  X"D0",  X"82",  X"96",  X"92",  X"94",  X"82",  X"7F",
  X"9E",  X"01",  X"9D",  X"80",  X"02",  X"A0",  X"80",  X"02",
  X"E6",  X"D4",  X"A2",  X"E8",  X"EA",  X"90",  X"92",  X"96",
  X"7F",  X"A4",  X"80",  X"02",  X"B0",  X"82",  X"80",  X"2A",
  X"EA",  X"80",  X"3A",  X"EA",  X"80",  X"02",  X"B0",  X"80",
  X"04",  X"82",  X"C4",  X"C4",  X"82",  X"80",  X"32",  X"C4",
  X"A4",  X"C2",  X"82",  X"C2",  X"C2",  X"80",  X"02",  X"80",
  X"1A",  X"A6",  X"D4",  X"E8",  X"EA",  X"90",  X"92",  X"7F",
  X"96",  X"80",  X"12",  X"82",  X"82",  X"C2",  X"C0",  X"81",
  X"91",  X"E8",  X"81",  X"81",  X"B0",  X"81",  X"81",  X"80",
  X"32",  X"C0",  X"C0",  X"81",  X"91",  X"E6",  X"10",  X"B6",
  X"03",  X"86",  X"84",  X"D0",  X"82",  X"98",  X"92",  X"94",
  X"96",  X"82",  X"7F",  X"9E",  X"01",  X"9D",  X"21",  X"40",
  X"90",  X"80",  X"08",  X"90",  X"13",  X"40",  X"92",  X"80",
  X"12",  X"80",  X"02",  X"80",  X"24",  X"F4",  X"82",  X"80",
  X"18",  X"82",  X"B4",  X"82",  X"B5",  X"B4",  X"C2",  X"F4",
  X"81",  X"91",  X"90",  X"13",  X"40",  X"92",  X"80",  X"12",
  X"80",  X"02",  X"83",  X"84",  X"12",  X"86",  X"F4",  X"81",
  X"91",  X"80",  X"32",  X"F4",  X"81",  X"91",  X"84",  X"03",
  X"82",  X"80",  X"08",  X"05",  X"03",  X"84",  X"82",  X"80",
  X"18",  X"88",  X"87",  X"88",  X"86",  X"85",  X"86",  X"84",
  X"82",  X"84",  X"83",  X"82",  X"C8",  X"C6",  X"C4",  X"C2",
  X"81",  X"91",  X"05",  X"03",  X"84",  X"82",  X"80",  X"18",
  X"9A",  X"89",  X"9A",  X"88",  X"87",  X"88",  X"86",  X"85",
  X"86",  X"84",  X"82",  X"84",  X"83",  X"82",  X"DA",  X"C8",
  X"C6",  X"C4",  X"C2",  X"81",  X"91",  X"86",  X"80",  X"38",
  X"82",  X"82",  X"82",  X"80",  X"08",  X"82",  X"86",  X"86",
  X"80",  X"38",  X"B0",  X"C2",  X"C4",  X"81",  X"91",  X"90",
  X"13",  X"40",  X"92",  X"80",  X"12",  X"80",  X"02",  X"83",
  X"80",  X"22",  X"F4",  X"84",  X"84",  X"80",  X"08",  X"84",
  X"81",  X"91",  X"90",  X"13",  X"40",  X"92",  X"80",  X"12",
  X"80",  X"02",  X"B0",  X"83",  X"86",  X"12",  X"84",  X"C2",
  X"80",  X"02",  X"82",  X"C0",  X"C2",  X"82",  X"B0",  X"C2",
  X"82",  X"C2",  X"B2",  X"C4",  X"81",  X"81",  X"03",  X"82",
  X"80",  X"08",  X"86",  X"85",  X"86",  X"84",  X"82",  X"84",
  X"83",  X"82",  X"C6",  X"C4",  X"C2",  X"81",  X"91",  X"82",
  X"80",  X"08",  X"82",  X"81",  X"91",  X"98",  X"9B",  X"98",
  X"9A",  X"89",  X"9A",  X"88",  X"87",  X"88",  X"86",  X"85",
  X"86",  X"84",  X"82",  X"84",  X"83",  X"82",  X"D8",  X"DA",
  X"C8",  X"C6",  X"C4",  X"C2",  X"81",  X"91",  X"82",  X"82",
  X"80",  X"18",  X"B0",  X"82",  X"82",  X"80",  X"18",  X"01",
  X"C2",  X"80",  X"12",  X"B0",  X"82",  X"C2",  X"82",  X"C2",
  X"82",  X"B0",  X"C2",  X"82",  X"C2",  X"B2",  X"C4",  X"C6",
  X"81",  X"81",  X"84",  X"80",  X"38",  X"B0",  X"F4",  X"C2",
  X"81",  X"91",  X"9D",  X"23",  X"D0",  X"80",  X"02",  X"A0",
  X"C2",  X"80",  X"02",  X"01",  X"C2",  X"85",  X"85",  X"80",
  X"02",  X"86",  X"C4",  X"80",  X"02",  X"01",  X"C2",  X"80",
  X"12",  X"80",  X"02",  X"82",  X"C2",  X"B0",  X"81",  X"81",
  X"C2",  X"C2",  X"81",  X"91",  X"C2",  X"82",  X"C0",  X"C2",
  X"81",  X"91",  X"40",  X"01",  X"10",  X"C2",  X"40",  X"90",
  X"10",  X"C2",  X"80",  X"02",  X"B0",  X"80",  X"32",  X"D2",
  X"86",  X"C4",  X"10",  X"C6",  X"80",  X"02",  X"86",  X"84",
  X"80",  X"22",  X"C0",  X"40",  X"D0",  X"C2",  X"C0",  X"86",
  X"C4",  X"C0",  X"C6",  X"86",  X"C4",  X"10",  X"C6",  X"9D",
  X"C2",  X"E6",  X"A0",  X"80",  X"14",  X"B0",  X"BA",  X"BB",
  X"82",  X"BA",  X"F4",  X"D2",  X"92",  X"90",  X"40",  X"A6",
  X"BA",  X"B0",  X"A2",  X"02",  X"B8",  X"2B",  X"A8",  X"AA",
  X"A4",  X"AC",  X"B6",  X"EE",  X"92",  X"40",  X"90",  X"93",
  X"AC",  X"40",  X"90",  X"C2",  X"87",  X"82",  X"B6",  X"84",
  X"AD",  X"84",  X"AC",  X"83",  X"88",  X"86",  X"B6",  X"C4",
  X"A8",  X"F6",  X"80",  X"A4",  X"AD",  X"1A",  X"B7",  X"80",
  X"12",  X"92",  X"84",  X"85",  X"82",  X"80",  X"3A",  X"E6",
  X"C4",  X"80",  X"02",  X"82",  X"10",  X"E6",  X"C4",  X"80",
  X"12",  X"82",  X"80",  X"0A",  X"A6",  X"E6",  X"92",  X"40",
  X"90",  X"80",  X"06",  X"17",  X"B0",  X"96",  X"82",  X"98",
  X"C8",  X"DA",  X"87",  X"85",  X"88",  X"84",  X"86",  X"86",
  X"86",  X"89",  X"84",  X"C6",  X"A2",  X"C4",  X"80",  X"82",
  X"1A",  X"99",  X"84",  X"85",  X"82",  X"C6",  X"80",  X"12",
  X"80",  X"3A",  X"E6",  X"C4",  X"80",  X"22",  X"82",  X"E6",
  X"81",  X"81",  X"C4",  X"80",  X"32",  X"E6",  X"82",  X"80",
  X"0A",  X"A6",  X"E6",  X"81",  X"81",  X"9D",  X"C2",  X"F2",
  X"F4",  X"80",  X"E2",  X"E0",  X"02",  X"D1",  X"C4",  X"C4",
  X"86",  X"D1",  X"C4",  X"85",  X"C4",  X"D3",  X"92",  X"40",
  X"90",  X"D3",  X"C0",  X"D1",  X"D1",  X"E4",  X"80",  X"06",
  X"82",  X"C0",  X"03",  X"84",  X"80",  X"02",  X"23",  X"95",
  X"D9",  X"97",  X"81",  X"01",  X"03",  X"82",  X"C2",  X"31",
  X"80",  X"02",  X"B0",  X"31",  X"B0",  X"F0",  X"81",  X"91",
  X"84",  X"C4",  X"E6",  X"90",  X"40",  X"92",  X"C0",  X"80",
  X"B0",  X"C4",  X"82",  X"02",  X"C2",  X"E4",  X"81",  X"81",
  X"D3",  X"03",  X"82",  X"C2",  X"C4",  X"80",  X"02",  X"03",
  X"31",  X"B0",  X"80",  X"02",  X"01",  X"C2",  X"80",  X"02",
  X"82",  X"82",  X"C2",  X"81",  X"81",  X"C2",  X"03",  X"A4",
  X"E4",  X"10",  X"D1",  X"D5",  X"D1",  X"D3",  X"D1",  X"D3",
  X"90",  X"96",  X"D8",  X"92",  X"94",  X"40",  X"98",  X"89",
  X"A8",  X"88",  X"D1",  X"D3",  X"D5",  X"12",  X"D7",  X"D3",
  X"C2",  X"C6",  X"86",  X"88",  X"84",  X"80",  X"DA",  X"04",
  X"85",  X"86",  X"84",  X"87",  X"85",  X"84",  X"C4",  X"80",
  X"DD",  X"06",  X"99",  X"D9",  X"88",  X"D8",  X"86",  X"1B",
  X"84",  X"84",  X"9A",  X"DA",  X"C4",  X"C8",  X"1B",  X"DD",
  X"05",  X"D9",  X"9D",  X"D9",  X"9D",  X"DB",  X"A1",  X"05",
  X"D9",  X"9D",  X"05",  X"D9",  X"99",  X"99",  X"DD",  X"81",
  X"9D",  X"DD",  X"01",  X"19",  X"E6",  X"9D",  X"81",  X"01",
  X"23",  X"A6",  X"84",  X"80",  X"18",  X"C4",  X"85",  X"07",
  X"86",  X"D9",  X"81",  X"01",  X"19",  X"C0",  X"A6",  X"82",
  X"B4",  X"82",  X"80",  X"06",  X"B2",  X"B4",  X"B2",  X"80",
  X"06",  X"86",  X"E6",  X"C0",  X"B4",  X"80",  X"18",  X"86",
  X"80",  X"04",  X"A4",  X"B6",  X"A4",  X"80",  X"02",  X"AE",
  X"04",  X"80",  X"80",  X"02",  X"80",  X"12",  X"88",  X"AE",
  X"9A",  X"88",  X"AC",  X"04",  X"DA",  X"C0",  X"80",  X"84",
  X"08",  X"82",  X"92",  X"83",  X"86",  X"80",  X"08",  X"84",
  X"80",  X"D2",  X"82",  X"D1",  X"A4",  X"D3",  X"D5",  X"D7",
  X"40",  X"90",  X"D0",  X"AA",  X"80",  X"D1",  X"D3",  X"D5",
  X"12",  X"D7",  X"80",  X"14",  X"C2",  X"80",  X"06",  X"05",
  X"83",  X"80",  X"84",  X"04",  X"D9",  X"95",  X"80",  X"A4",
  X"95",  X"D5",  X"9D",  X"9D",  X"91",  X"D8",  X"82",  X"02",
  X"C2",  X"1B",  X"D5",  X"91",  X"D5",  X"81",  X"01",  X"13",
  X"82",  X"86",  X"10",  X"A2",  X"D5",  X"91",  X"D5",  X"81",
  X"01",  X"33",  X"E6",  X"95",  X"82",  X"80",  X"95",  X"D5",
  X"9D",  X"9D",  X"91",  X"C8",  X"84",  X"C4",  X"12",  X"A4",
  X"91",  X"81",  X"01",  X"29",  X"C2",  X"81",  X"01",  X"23",
  X"E6",  X"D5",  X"DA",  X"80",  X"32",  X"C2",  X"10",  X"E6",
  X"31",  X"80",  X"02",  X"B0",  X"10",  X"31",  X"D5",  X"03",
  X"88",  X"C0",  X"D8",  X"84",  X"86",  X"1B",  X"9A",  X"84",
  X"10",  X"C2",  X"C6",  X"A4",  X"B6",  X"AE",  X"AC",  X"B8",
  X"C0",  X"92",  X"D1",  X"D3",  X"D5",  X"D7",  X"40",  X"90",
  X"D0",  X"AA",  X"80",  X"D1",  X"D3",  X"D5",  X"02",  X"D7",
  X"80",  X"04",  X"82",  X"83",  X"05",  X"99",  X"84",  X"9B",
  X"D1",  X"83",  X"80",  X"12",  X"86",  X"80",  X"22",  X"91",
  X"05",  X"84",  X"80",  X"02",  X"83",  X"DD",  X"91",  X"86",
  X"80",  X"12",  X"84",  X"91",  X"C2",  X"80",  X"22",  X"C6",
  X"03",  X"D9",  X"81",  X"01",  X"19",  X"01",  X"80",  X"04",
  X"C4",  X"80",  X"04",  X"86",  X"C6",  X"1B",  X"D9",  X"91",
  X"03",  X"D9",  X"9D",  X"9D",  X"D9",  X"A1",  X"E1",  X"03",
  X"D8",  X"98",  X"82",  X"10",  X"C2",  X"C6",  X"03",  X"80",
  X"D9",  X"9D",  X"9D",  X"D9",  X"A1",  X"E1",  X"03",  X"D8",
  X"12",  X"98",  X"D8",  X"03",  X"D9",  X"91",  X"D9",  X"81",
  X"01",  X"2D",  X"C0",  X"99",  X"81",  X"01",  X"19",  X"01",
  X"C0",  X"A2",  X"A6",  X"EE",  X"A4",  X"10",  X"B8",  X"80",
  X"12",  X"80",  X"E2",  X"F2",  X"C0",  X"80",  X"04",  X"D8",
  X"80",  X"04",  X"80",  X"04",  X"82",  X"82",  X"DA",  X"9A",
  X"DA",  X"B4",  X"B2",  X"C2",  X"80",  X"04",  X"80",  X"02",
  X"80",  X"04",  X"D2",  X"D1",  X"D3",  X"94",  X"40",  X"90",
  X"D0",  X"94",  X"90",  X"40",  X"D2",  X"92",  X"A4",  X"40",
  X"90",  X"D3",  X"D1",  X"A8",  X"C4",  X"94",  X"12",  X"92",
  X"D1",  X"D3",  X"90",  X"40",  X"92",  X"C6",  X"A2",  X"80",
  X"D1",  X"04",  X"D3",  X"92",  X"94",  X"40",  X"90",  X"D3",
  X"D1",  X"A2",  X"80",  X"24",  X"D3",  X"C0",  X"DA",  X"80",
  X"12",  X"82",  X"82",  X"82",  X"12",  X"84",  X"C6",  X"86",
  X"C6",  X"B4",  X"B2",  X"80",  X"04",  X"92",  X"D1",  X"D3",
  X"94",  X"40",  X"90",  X"D3",  X"D1",  X"A8",  X"80",  X"04",
  X"92",  X"D1",  X"D3",  X"94",  X"40",  X"90",  X"D3",  X"D1",
  X"A2",  X"C8",  X"80",  X"32",  X"D1",  X"80",  X"04",  X"80",
  X"80",  X"A4",  X"02",  X"AE",  X"D8",  X"80",  X"04",  X"D2",
  X"D1",  X"D3",  X"94",  X"40",  X"90",  X"D3",  X"D0",  X"D1",
  X"DA",  X"80",  X"12",  X"EE",  X"D3",  X"F8",  X"A4",  X"B4",
  X"C6",  X"B2",  X"92",  X"7F",  X"90",  X"90",  X"92",  X"D0",
  X"40",  X"90",  X"92",  X"D0",  X"94",  X"40",  X"90",  X"C4",
  X"80",  X"82",  X"02",  X"84",  X"C4",  X"92",  X"40",  X"90",
  X"C4",  X"80",  X"12",  X"DA",  X"80",  X"12",  X"80",  X"80",
  X"02",  X"C8",  X"80",  X"06",  X"80",  X"12",  X"80",  X"80",
  X"12",  X"80",  X"80",  X"02",  X"80",  X"14",  X"DA",  X"80",
  X"DA",  X"02",  X"A4",  X"92",  X"90",  X"94",  X"40",  X"96",
  X"80",  X"02",  X"A8",  X"92",  X"94",  X"96",  X"40",  X"90",
  X"92",  X"B8",  X"94",  X"90",  X"96",  X"40",  X"B4",  X"10",
  X"AE",  X"B2",  X"C6",  X"10",  X"C0",  X"05",  X"D9",  X"99",
  X"82",  X"10",  X"86",  X"02",  X"88",  X"A4",  X"AE",  X"C8",
  X"AC",  X"10",  X"B8",  X"90",  X"94",  X"96",  X"40",  X"AE",
  X"A8",  X"92",  X"7F",  X"90",  X"90",  X"D0",  X"80",  X"D0",
  X"92",  X"06",  X"A4",  X"EE",  X"B8",  X"92",  X"94",  X"40",
  X"90",  X"92",  X"40",  X"A8",  X"80",  X"34",  X"C2",  X"30",
  X"C2",  X"80",  X"C4",  X"12",  X"82",  X"80",  X"32",  X"A4",
  X"82",  X"C2",  X"A6",  X"92",  X"40",  X"90",  X"80",  X"02",
  X"80",  X"02",  X"80",  X"02",  X"92",  X"40",  X"90",  X"92",
  X"E6",  X"40",  X"90",  X"10",  X"90",  X"04",  X"DA",  X"82",
  X"80",  X"16",  X"A2",  X"C6",  X"82",  X"84",  X"86",  X"C4",
  X"C6",  X"A2",  X"88",  X"C8",  X"80",  X"06",  X"82",  X"F2",
  X"82",  X"D1",  X"D3",  X"B4",  X"B2",  X"90",  X"40",  X"92",
  X"D3",  X"D0",  X"10",  X"D1",  X"E6",  X"84",  X"80",  X"22",
  X"99",  X"82",  X"83",  X"07",  X"86",  X"D9",  X"03",  X"DD",
  X"9D",  X"99",  X"D9",  X"99",  X"99",  X"C6",  X"82",  X"C2",
  X"D8",  X"D1",  X"91",  X"81",  X"01",  X"0D",  X"A4",  X"09",
  X"DD",  X"9D",  X"81",  X"01",  X"0D",  X"80",  X"04",  X"1B",
  X"88",  X"E1",  X"10",  X"82",  X"DD",  X"9D",  X"81",  X"01",
  X"29",  X"E6",  X"36",  X"91",  X"99",  X"9D",  X"DD",  X"9D",
  X"99",  X"91",  X"82",  X"81",  X"80",  X"D8",  X"86",  X"C6",
  X"01",  X"19",  X"A4",  X"10",  X"90",  X"C8",  X"80",  X"32",
  X"C0",  X"D1",  X"05",  X"C2",  X"80",  X"32",  X"C0",  X"05",
  X"80",  X"22",  X"C0",  X"98",  X"B2",  X"B4",  X"10",  X"D8",
  X"C2",  X"80",  X"C4",  X"12",  X"82",  X"80",  X"32",  X"A4",
  X"82",  X"A6",  X"C2",  X"84",  X"10",  X"82",  X"91",  X"10",
  X"93",  X"92",  X"C2",  X"40",  X"90",  X"C2",  X"10",  X"84",
  X"80",  X"36",  X"95",  X"80",  X"12",  X"03",  X"D5",  X"99",
  X"81",  X"01",  X"17",  X"C0",  X"A2",  X"EE",  X"82",  X"A6",
  X"C2",  X"A4",  X"10",  X"B8",  X"84",  X"82",  X"80",  X"04",
  X"C4",  X"82",  X"84",  X"B4",  X"B2",  X"10",  X"C4",  X"92",
  X"90",  X"94",  X"96",  X"40",  X"B4",  X"B8",  X"10",  X"AE",
  X"91",  X"93",  X"82",  X"02",  X"86",  X"84",  X"07",  X"85",
  X"86",  X"D1",  X"83",  X"91",  X"80",  X"02",  X"86",  X"05",
  X"84",  X"80",  X"02",  X"83",  X"D9",  X"91",  X"86",  X"80",
  X"12",  X"84",  X"10",  X"C2",  X"D9",  X"99",  X"91",  X"80",
  X"A4",  X"C6",  X"82",  X"07",  X"86",  X"C2",  X"D8",  X"82",
  X"83",  X"E1",  X"DD",  X"02",  X"A1",  X"1B",  X"DD",  X"82",
  X"91",  X"99",  X"D9",  X"99",  X"C8",  X"86",  X"C6",  X"82",
  X"80",  X"12",  X"91",  X"82",  X"A4",  X"03",  X"D9",  X"9D",
  X"81",  X"01",  X"2D",  X"E6",  X"99",  X"81",  X"01",  X"19",
  X"01",  X"10",  X"C2",  X"A4",  X"C2",  X"80",  X"02",  X"82",
  X"10",  X"90",  X"05",  X"DD",  X"10",  X"99",  X"AE",  X"80",
  X"04",  X"88",  X"F8",  X"10",  X"AC",  X"10",  X"AE",  X"10",
  X"E6",  X"C2",  X"82",  X"83",  X"82",  X"D0",  X"D1",  X"40",
  X"D3",  X"82",  X"D3",  X"82",  X"10",  X"D1",  X"D3",  X"90",
  X"40",  X"92",  X"D1",  X"80",  X"16",  X"D3",  X"92",  X"90",
  X"94",  X"40",  X"96",  X"A6",  X"A8",  X"80",  X"EC",  X"D1",
  X"02",  X"D3",  X"D2",  X"90",  X"94",  X"40",  X"96",  X"D3",
  X"D0",  X"10",  X"D1",  X"80",  X"82",  X"10",  X"A4",  X"98",
  X"AC",  X"D8",  X"10",  X"B8",  X"D4",  X"92",  X"D1",  X"D3",
  X"40",  X"90",  X"D3",  X"A8",  X"10",  X"D1",  X"04",  X"80",
  X"80",  X"12",  X"92",  X"94",  X"96",  X"40",  X"90",  X"A2",
  X"90",  X"40",  X"92",  X"80",  X"34",  X"EE",  X"10",  X"A6",
  X"D1",  X"D3",  X"40",  X"90",  X"D1",  X"A8",  X"10",  X"D3",
  X"D8",  X"80",  X"22",  X"C2",  X"82",  X"E2",  X"10",  X"F2",
  X"80",  X"04",  X"92",  X"94",  X"40",  X"90",  X"92",  X"40",
  X"A8",  X"80",  X"04",  X"C4",  X"80",  X"02",  X"84",  X"C4",
  X"C6",  X"C6",  X"10",  X"A4",  X"32",  X"C2",  X"C2",  X"80",
  X"12",  X"C2",  X"10",  X"80",  X"A4",  X"C2",  X"80",  X"02",
  X"82",  X"10",  X"92",  X"84",  X"10",  X"C4",  X"D2",  X"D3",
  X"D1",  X"40",  X"90",  X"C4",  X"D4",  X"92",  X"A4",  X"94",
  X"90",  X"40",  X"95",  X"90",  X"92",  X"40",  X"94",  X"D3",
  X"10",  X"AE",  X"84",  X"E2",  X"82",  X"10",  X"F2",  X"C8",
  X"80",  X"02",  X"D8",  X"82",  X"C2",  X"10",  X"A4",  X"82",
  X"C2",  X"10",  X"A4",  X"80",  X"02",  X"D8",  X"83",  X"82",
  X"83",  X"88",  X"C8",  X"10",  X"A4",  X"12",  X"C6",  X"C2",
  X"80",  X"22",  X"C6",  X"10",  X"C4",  X"80",  X"92",  X"82",
  X"10",  X"A4",  X"02",  X"80",  X"10",  X"84",  X"9D",  X"80",
  X"02",  X"03",  X"C2",  X"80",  X"02",  X"01",  X"03",  X"D0",
  X"80",  X"22",  X"C6",  X"C2",  X"80",  X"02",  X"01",  X"C6",
  X"83",  X"85",  X"80",  X"22",  X"83",  X"E2",  X"80",  X"02",
  X"80",  X"E0",  X"E2",  X"A0",  X"12",  X"82",  X"C2",  X"80",
  X"14",  X"C2",  X"10",  X"80",  X"A0",  X"80",  X"24",  X"C6",
  X"C2",  X"D0",  X"92",  X"9F",  X"94",  X"80",  X"14",  X"A2",
  X"C4",  X"84",  X"82",  X"80",  X"12",  X"C4",  X"40",  X"90",
  X"10",  X"82",  X"83",  X"80",  X"02",  X"82",  X"81",  X"91",
  X"80",  X"12",  X"82",  X"40",  X"90",  X"82",  X"81",  X"91",
  X"40",  X"90",  X"10",  X"03",  X"40",  X"01",  X"10",  X"C6",
  X"F0",  X"03",  X"40",  X"93",  X"01",  X"13",  X"92",  X"82",
  X"40",  X"9E",  X"01",  X"03",  X"D0",  X"82",  X"7F",  X"9E",
  X"01",  X"9D",  X"C2",  X"80",  X"12",  X"01",  X"40",  X"90",
  X"81",  X"91",  X"11",  X"90",  X"82",  X"40",  X"9E",  X"01",
  X"9D",  X"03",  X"D0",  X"13",  X"40",  X"92",  X"7F",  X"81",
  X"01",  X"9D",  X"C2",  X"80",  X"12",  X"01",  X"40",  X"90",
  X"81",  X"91",  X"11",  X"90",  X"82",  X"40",  X"9E",  X"01",
  X"9D",  X"7F",  X"33",  X"03",  X"F0",  X"40",  X"93",  X"01",
  X"9D",  X"03",  X"82",  X"C2",  X"03",  X"82",  X"C2",  X"03",
  X"82",  X"F0",  X"C2",  X"F2",  X"F4",  X"C0",  X"C0",  X"C0",
  X"C0",  X"C0",  X"C0",  X"03",  X"82",  X"C2",  X"A0",  X"40",
  X"90",  X"90",  X"40",  X"92",  X"92",  X"40",  X"90",  X"40",
  X"90",  X"81",  X"81",  X"9D",  X"03",  X"82",  X"C2",  X"82",
  X"C2",  X"82",  X"D0",  X"C2",  X"C0",  X"82",  X"C2",  X"96",
  X"92",  X"7F",  X"94",  X"D0",  X"96",  X"B6",  X"92",  X"7F",
  X"94",  X"F0",  X"B2",  X"7F",  X"95",  X"01",  X"9D",  X"83",
  X"A1",  X"A0",  X"83",  X"90",  X"A0",  X"7F",  X"92",  X"B0",
  X"02",  X"90",  X"F2",  X"C0",  X"D0",  X"94",  X"40",  X"92",
  X"81",  X"81",  X"9D",  X"7F",  X"01",  X"03",  X"E2",  X"C2",
  X"80",  X"02",  X"01",  X"A2",  X"C2",  X"82",  X"1C",  X"E0",
  X"10",  X"D0",  X"0C",  X"A0",  X"C4",  X"80",  X"12",  X"82",
  X"82",  X"C2",  X"82",  X"C2",  X"A2",  X"40",  X"90",  X"92",
  X"40",  X"90",  X"92",  X"40",  X"90",  X"40",  X"90",  X"7F",
  X"01",  X"C0",  X"C0",  X"C0",  X"C0",  X"C0",  X"C0",  X"C0",
  X"C0",  X"C0",  X"C0",  X"81",  X"91",  X"D0",  X"80",  X"22",
  X"90",  X"10",  X"A2",  X"7F",  X"90",  X"10",  X"A2",  X"7F",
  X"92",  X"80",  X"12",  X"D0",  X"7F",  X"A0",  X"82",  X"10",
  X"C2",  X"9D",  X"7F",  X"90",  X"21",  X"A0",  X"C2",  X"E2",
  X"A2",  X"82",  X"B2",  X"B2",  X"B2",  X"80",  X"04",  X"90",
  X"7F",  X"92",  X"C2",  X"82",  X"80",  X"02",  X"90",  X"90",
  X"7F",  X"B0",  X"81",  X"81",  X"7F",  X"92",  X"80",  X"02",
  X"A2",  X"C4",  X"A2",  X"03",  X"E2",  X"90",  X"B0",  X"C4",
  X"B2",  X"7F",  X"F2",  X"81",  X"81",  X"90",  X"7F",  X"92",
  X"C2",  X"84",  X"80",  X"04",  X"07",  X"C6",  X"90",  X"07",
  X"84",  X"D0",  X"10",  X"C4",  X"9D",  X"80",  X"02",  X"01",
  X"7F",  X"90",  X"84",  X"D8",  X"82",  X"09",  X"86",  X"88",
  X"DA",  X"D6",  X"80",  X"02",  X"9A",  X"DA",  X"80",  X"12",
  X"98",  X"D8",  X"84",  X"82",  X"D6",  X"98",  X"80",  X"02",
  X"98",  X"D4",  X"D4",  X"98",  X"D6",  X"96",  X"D6",  X"80",
  X"32",  X"86",  X"80",  X"02",  X"82",  X"DA",  X"C6",  X"C6",
  X"DA",  X"86",  X"C2",  X"80",  X"12",  X"C6",  X"80",  X"28",
  X"83",  X"87",  X"80",  X"18",  X"98",  X"99",  X"98",  X"9B",
  X"9A",  X"C6",  X"80",  X"32",  X"C8",  X"10",  X"DA",  X"80",
  X"22",  X"C2",  X"C8",  X"88",  X"80",  X"2A",  X"C6",  X"C2",
  X"C2",  X"C6",  X"C4",  X"C4",  X"7F",  X"81",  X"81",  X"81",
  X"DA",  X"17",  X"96",  X"80",  X"32",  X"C6",  X"C4",  X"C4",
  X"C2",  X"DA",  X"82",  X"DA",  X"C2",  X"7F",  X"81",  X"87",
  X"86",  X"DA",  X"C6",  X"DA",  X"D8",  X"C4",  X"C4",  X"83",
  X"84",  X"83",  X"82",  X"C2",  X"7F",  X"81",  X"80",  X"12",
  X"82",  X"D8",  X"84",  X"DA",  X"C6",  X"82",  X"C6",  X"DA",
  X"C4",  X"86",  X"C6",  X"05",  X"C4",  X"80",  X"0A",  X"03",
  X"D2",  X"7F",  X"90",  X"7F",  X"81",  X"80",  X"08",  X"9B",
  X"80",  X"18",  X"80",  X"99",  X"98",  X"10",  X"9B",  X"99",
  X"82",  X"83",  X"82",  X"C2",  X"10",  X"82",  X"18",  X"80",
  X"99",  X"98",  X"10",  X"9B",  X"9A",  X"18",  X"98",  X"99",
  X"98",  X"10",  X"9B",  X"9D",  X"C2",  X"80",  X"02",  X"A0",
  X"C4",  X"80",  X"02",  X"82",  X"C6",  X"80",  X"02",  X"90",
  X"80",  X"E2",  X"A6",  X"02",  X"A4",  X"80",  X"02",  X"92",
  X"80",  X"08",  X"94",  X"94",  X"C2",  X"9F",  X"D0",  X"80",
  X"04",  X"A4",  X"C2",  X"82",  X"80",  X"02",  X"C2",  X"A6",
  X"80",  X"12",  X"92",  X"E6",  X"E4",  X"10",  X"A2",  X"B0",
  X"81",  X"81",  X"2D",  X"80",  X"AC",  X"02",  X"A8",  X"AE",
  X"AC",  X"A6",  X"80",  X"22",  X"EC",  X"80",  X"02",  X"90",
  X"80",  X"08",  X"AA",  X"AA",  X"D4",  X"E4",  X"A4",  X"80",
  X"04",  X"D0",  X"C2",  X"80",  X"08",  X"80",  X"92",  X"40",
  X"94",  X"C2",  X"82",  X"C2",  X"7F",  X"90",  X"80",  X"32",
  X"C2",  X"A8",  X"02",  X"01",  X"C2",  X"82",  X"80",  X"02",
  X"C2",  X"A6",  X"80",  X"12",  X"AC",  X"EC",  X"E6",  X"AE",
  X"10",  X"A2",  X"D0",  X"80",  X"1A",  X"94",  X"AA",  X"A6",
  X"94",  X"40",  X"92",  X"C4",  X"C2",  X"A6",  X"AA",  X"E6",
  X"EA",  X"A6",  X"AA",  X"C2",  X"A6",  X"80",  X"02",  X"E6",
  X"C2",  X"A4",  X"A8",  X"80",  X"22",  X"E8",  X"83",  X"83",
  X"80",  X"02",  X"E6",  X"80",  X"08",  X"AA",  X"80",  X"22",
  X"D0",  X"D2",  X"EA",  X"D0",  X"AA",  X"A6",  X"40",  X"94",
  X"82",  X"02",  X"90",  X"E6",  X"C2",  X"D0",  X"E4",  X"A6",
  X"10",  X"AA",  X"E4",  X"10",  X"A2",  X"80",  X"D0",  X"1A",
  X"AA",  X"C2",  X"80",  X"28",  X"D4",  X"92",  X"40",  X"94",
  X"C2",  X"82",  X"C2",  X"7F",  X"90",  X"80",  X"22",  X"C2",
  X"C2",  X"82",  X"C2",  X"81",  X"91",  X"D4",  X"80",  X"0A",
  X"92",  X"C2",  X"D0",  X"9F",  X"92",  X"A6",  X"24",  X"C2",
  X"10",  X"AA",  X"40",  X"94",  X"C4",  X"C2",  X"84",  X"82",
  X"C4",  X"C2",  X"A6",  X"10",  X"AA",  X"80",  X"06",  X"92",
  X"C2",  X"D0",  X"9F",  X"92",  X"A4",  X"24",  X"C2",  X"A8",
  X"32",  X"C2",  X"7F",  X"90",  X"80",  X"12",  X"AE",  X"10",
  X"C2",  X"40",  X"94",  X"C4",  X"C2",  X"84",  X"82",  X"C4",
  X"C2",  X"10",  X"A4",  X"92",  X"94",  X"40",  X"A8",  X"80",
  X"02",  X"AE",  X"A8",  X"10",  X"A8",  X"90",  X"7F",  X"B0",
  X"80",  X"12",  X"01",  X"C2",  X"10",  X"84",  X"D0",  X"7F",
  X"D2",  X"10",  X"C2",  X"9D",  X"7F",  X"A0",  X"A6",  X"02",
  X"B0",  X"E4",  X"A4",  X"1C",  X"E2",  X"10",  X"E6",  X"C4",
  X"92",  X"80",  X"02",  X"90",  X"9F",  X"01",  X"C2",  X"B0",
  X"80",  X"02",  X"A8",  X"A4",  X"2C",  X"E6",  X"A2",  X"C2",
  X"85",  X"80",  X"22",  X"A4",  X"85",  X"80",  X"32",  X"C4",
  X"A8",  X"40",  X"90",  X"C2",  X"80",  X"12",  X"C2",  X"40",
  X"90",  X"A4",  X"3C",  X"A2",  X"E6",  X"80",  X"32",  X"E4",
  X"7F",  X"01",  X"81",  X"81",  X"9D",  X"7F",  X"01",  X"A4",
  X"02",  X"B0",  X"E2",  X"A2",  X"1C",  X"E0",  X"10",  X"E4",
  X"C4",  X"80",  X"02",  X"90",  X"9F",  X"01",  X"C2",  X"B0",
  X"80",  X"02",  X"A6",  X"A2",  X"2C",  X"E4",  X"A0",  X"C2",
  X"85",  X"80",  X"22",  X"A2",  X"85",  X"80",  X"32",  X"C4",
  X"A6",  X"40",  X"90",  X"C2",  X"80",  X"12",  X"C2",  X"40",
  X"90",  X"A2",  X"3C",  X"A0",  X"E4",  X"80",  X"32",  X"E2",
  X"7F",  X"01",  X"81",  X"81",  X"03",  X"81",  X"D0",  X"11",
  X"81",  X"90",  X"11",  X"81",  X"90",  X"9D",  X"A0",  X"80",
  X"31",  X"02",  X"B0",  X"90",  X"92",  X"40",  X"23",  X"80",
  X"12",  X"90",  X"F4",  X"F2",  X"81",  X"91",  X"13",  X"B0",
  X"40",  X"92",  X"80",  X"22",  X"F4",  X"81",  X"81",  X"82",
  X"05",  X"D0",  X"94",  X"92",  X"82",  X"7F",  X"9E",  X"01",
  X"9D",  X"C2",  X"80",  X"32",  X"82",  X"D2",  X"80",  X"06",
  X"21",  X"D0",  X"40",  X"94",  X"80",  X"06",  X"C4",  X"03",
  X"82",  X"05",  X"84",  X"80",  X"05",  X"A2",  X"80",  X"22",
  X"C4",  X"C2",  X"82",  X"10",  X"C2",  X"C2",  X"82",  X"A2",
  X"C2",  X"D0",  X"7F",  X"92",  X"80",  X"02",  X"03",  X"C4",
  X"C2",  X"84",  X"D0",  X"D0",  X"C4",  X"05",  X"84",  X"C4",
  X"82",  X"80",  X"02",  X"C2",  X"40",  X"D0",  X"80",  X"02",
  X"01",  X"C2",  X"82",  X"C2",  X"81",  X"81",  X"C2",  X"C2",
  X"82",  X"C2",  X"81",  X"81",  X"03",  X"82",  X"80",  X"12",
  X"C2",  X"82",  X"84",  X"C4",  X"10",  X"C2",  X"C4",  X"84",
  X"82",  X"C2",  X"C2",  X"C4",  X"82",  X"C2",  X"81",  X"81",
  X"9D",  X"B2",  X"80",  X"08",  X"82",  X"80",  X"12",  X"9B",
  X"09",  X"9A",  X"07",  X"9B",  X"88",  X"9A",  X"86",  X"9B",
  X"9A",  X"C2",  X"82",  X"84",  X"82",  X"80",  X"02",  X"B4",
  X"C2",  X"80",  X"02",  X"01",  X"C2",  X"80",  X"02",  X"82",
  X"C2",  X"80",  X"02",  X"82",  X"C2",  X"80",  X"02",  X"82",
  X"80",  X"18",  X"B0",  X"82",  X"80",  X"32",  X"C4",  X"81",
  X"91",  X"80",  X"02",  X"82",  X"C4",  X"80",  X"12",  X"B4",
  X"81",  X"91",  X"81",  X"81",  X"9D",  X"80",  X"9A",  X"88",
  X"08",  X"86",  X"82",  X"80",  X"02",  X"84",  X"80",  X"02",
  X"82",  X"C4",  X"C4",  X"82",  X"80",  X"32",  X"C4",  X"81",
  X"81",  X"82",  X"DA",  X"DA",  X"86",  X"80",  X"DA",  X"DA",
  X"DA",  X"DA",  X"DA",  X"DA",  X"84",  X"18",  X"82",  X"B4",
  X"9B",  X"83",  X"9A",  X"B4",  X"9B",  X"80",  X"88",  X"86",
  X"08",  X"9A",  X"82",  X"C4",  X"C4",  X"82",  X"84",  X"80",
  X"38",  X"C4",  X"B4",  X"83",  X"87",  X"82",  X"86",  X"83",
  X"88",  X"10",  X"9A",  X"9D",  X"80",  X"9A",  X"88",  X"08",
  X"86",  X"82",  X"80",  X"1A",  X"80",  X"80",  X"02",  X"86",
  X"84",  X"82",  X"C8",  X"84",  X"86",  X"80",  X"12",  X"C8",
  X"81",  X"81",  X"80",  X"18",  X"82",  X"80",  X"02",  X"82",
  X"C4",  X"C4",  X"82",  X"80",  X"32",  X"C4",  X"81",  X"81",
  X"80",  X"12",  X"80",  X"86",  X"84",  X"82",  X"C8",  X"C8",
  X"86",  X"80",  X"C8",  X"C8",  X"C8",  X"C8",  X"C8",  X"C8",
  X"84",  X"18",  X"82",  X"B4",  X"9B",  X"83",  X"9A",  X"B4",
  X"9B",  X"80",  X"88",  X"86",  X"08",  X"9A",  X"82",  X"C4",
  X"C4",  X"82",  X"84",  X"80",  X"38",  X"C4",  X"B4",  X"83",
  X"87",  X"82",  X"86",  X"83",  X"88",  X"10",  X"9A",  X"9D",
  X"86",  X"80",  X"08",  X"84",  X"80",  X"32",  X"82",  X"83",
  X"82",  X"80",  X"85",  X"9A",  X"84",  X"88",  X"08",  X"82",
  X"C4",  X"C4",  X"C4",  X"C4",  X"88",  X"80",  X"18",  X"82",
  X"82",  X"B4",  X"9A",  X"80",  X"9A",  X"08",  X"9A",  X"82",
  X"C4",  X"82",  X"88",  X"80",  X"38",  X"C4",  X"82",  X"B4",
  X"82",  X"82",  X"9A",  X"84",  X"80",  X"02",  X"82",  X"C6",
  X"82",  X"80",  X"32",  X"C6",  X"81",  X"81",  X"80",  X"02",
  X"01",  X"C4",  X"C2",  X"83",  X"C6",  X"C6",  X"D2",  X"81",
  X"01",  X"82",  X"05",  X"80",  X"12",  X"90",  X"83",  X"90",
  X"05",  X"80",  X"12",  X"05",  X"90",  X"83",  X"80",  X"12",
  X"05",  X"90",  X"83",  X"80",  X"12",  X"80",  X"90",  X"83",
  X"80",  X"06",  X"05",  X"80",  X"02",  X"90",  X"81",  X"01",
  X"81",  X"90",  X"C2",  X"80",  X"02",  X"05",  X"80",  X"12",
  X"84",  X"80",  X"12",  X"84",  X"83",  X"C2",  X"81",  X"90",
  X"84",  X"80",  X"02",  X"84",  X"80",  X"12",  X"80",  X"84",
  X"83",  X"80",  X"12",  X"80",  X"84",  X"83",  X"80",  X"12",
  X"80",  X"84",  X"83",  X"80",  X"32",  X"C2",  X"83",  X"80",
  X"02",  X"84",  X"C2",  X"81",  X"90",  X"83",  X"80",  X"12",
  X"84",  X"10",  X"84",  X"84",  X"81",  X"90",  X"83",  X"84",
  X"C2",  X"81",  X"90",  X"9D",  X"82",  X"C4",  X"F0",  X"B0",
  X"12",  X"84",  X"85",  X"86",  X"84",  X"86",  X"84",  X"82",
  X"84",  X"86",  X"DA",  X"C8",  X"80",  X"12",  X"80",  X"0A",
  X"84",  X"81",  X"81",  X"80",  X"B0",  X"B0",  X"81",  X"81",
  X"03",  X"05",  X"82",  X"82",  X"80",  X"04",  X"9C",  X"84",
  X"86",  X"C4",  X"C1",  X"81",  X"9C",  X"82",  X"83",  X"80",
  X"04",  X"09",  X"82",  X"80",  X"04",  X"88",  X"84",  X"86",
  X"C4",  X"C1",  X"81",  X"9C",  X"82",  X"84",  X"89",  X"10",
  X"86",  X"86",  X"85",  X"C4",  X"C1",  X"81",  X"9C",  X"9D",
  X"E0",  X"A0",  X"A1",  X"E2",  X"7F",  X"90",  X"82",  X"82",
  X"C2",  X"A0",  X"80",  X"14",  X"B0",  X"84",  X"80",  X"84",
  X"1A",  X"82",  X"C2",  X"83",  X"9B",  X"90",  X"09",  X"A3",
  X"84",  X"86",  X"C4",  X"C1",  X"81",  X"81",  X"80",  X"0A",
  X"82",  X"90",  X"02",  X"09",  X"84",  X"80",  X"84",  X"08",
  X"88",  X"C8",  X"89",  X"9B",  X"83",  X"05",  X"91",  X"86",
  X"90",  X"84",  X"C4",  X"C1",  X"81",  X"81",  X"09",  X"86",
  X"84",  X"C4",  X"C1",  X"81",  X"81",  X"C2",  X"90",  X"02",
  X"A0",  X"10",  X"84",  X"9D",  X"92",  X"7F",  X"90",  X"91",
  X"92",  X"90",  X"C3",  X"7F",  X"D1",  X"C6",  X"C4",  X"C2",
  X"C8",  X"82",  X"84",  X"D1",  X"85",  X"D3",  X"82",  X"80",
  X"04",  X"99",  X"D1",  X"83",  X"C4",  X"82",  X"C2",  X"D5",
  X"91",  X"81",  X"81",  X"81",  X"D9",  X"83",  X"C4",  X"82",
  X"C2",  X"D9",  X"81",  X"81",  X"81",  X"81",  X"80",  X"04",
  X"03",  X"C1",  X"03",  X"D1",  X"90",  X"12",  X"81",  X"81",
  X"01",  X"91",  X"03",  X"82",  X"81",  X"C1",  X"9D",  X"C2",
  X"80",  X"02",  X"A0",  X"85",  X"F0",  X"80",  X"02",  X"90",
  X"C6",  X"C6",  X"C0",  X"C0",  X"81",  X"81",  X"90",  X"92",
  X"40",  X"94",  X"D0",  X"82",  X"80",  X"12",  X"B0",  X"81",
  X"81",  X"92",  X"A0",  X"A1",  X"94",  X"40",  X"95",  X"B0",
  X"02",  X"01",  X"F2",  X"E0",  X"C0",  X"C0",  X"81",  X"81",
  X"9D",  X"92",  X"90",  X"F2",  X"7F",  X"F4",  X"05",  X"84",
  X"C4",  X"07",  X"A2",  X"82",  X"A5",  X"80",  X"02",  X"B0",
  X"07",  X"84",  X"C4",  X"80",  X"02",  X"01",  X"E2",  X"7F",
  X"90",  X"80",  X"12",  X"C2",  X"C2",  X"C2",  X"C2",  X"80",
  X"C2",  X"A0",  X"A0",  X"80",  X"12",  X"E0",  X"90",  X"82",
  X"D0",  X"83",  X"82",  X"7F",  X"D0",  X"A1",  X"A0",  X"E0",
  X"81",  X"81",  X"7F",  X"90",  X"C2",  X"C2",  X"82",  X"C2",
  X"90",  X"80",  X"02",  X"A0",  X"A4",  X"A4",  X"E4",  X"82",
  X"90",  X"D0",  X"81",  X"81",  X"C6",  X"84",  X"85",  X"84",
  X"C4",  X"83",  X"10",  X"C2",  X"9D",  X"E2",  X"C2",  X"A2",
  X"02",  X"90",  X"80",  X"06",  X"82",  X"A2",  X"A0",  X"7F",
  X"D2",  X"C8",  X"D2",  X"82",  X"E2",  X"83",  X"92",  X"B2",
  X"93",  X"19",  X"92",  X"B2",  X"92",  X"98",  X"B4",  X"82",
  X"84",  X"DA",  X"C6",  X"97",  X"9A",  X"95",  X"86",  X"96",
  X"86",  X"86",  X"9B",  X"84",  X"C6",  X"B4",  X"C4",  X"A0",
  X"82",  X"80",  X"18",  X"85",  X"80",  X"3A",  X"C4",  X"19",
  X"98",  X"C6",  X"9B",  X"86",  X"86",  X"85",  X"84",  X"C6",
  X"A0",  X"C4",  X"80",  X"82",  X"18",  X"85",  X"C4",  X"80",
  X"12",  X"82",  X"82",  X"C4",  X"80",  X"02",  X"88",  X"C8",
  X"81",  X"91",  X"82",  X"A0",  X"83",  X"84",  X"82",  X"84",
  X"82",  X"82",  X"84",  X"C8",  X"C6",  X"80",  X"12",  X"80",
  X"0A",  X"82",  X"7F",  X"92",  X"82",  X"C0",  X"C2",  X"81",
  X"91",  X"80",  X"1A",  X"82",  X"A2",  X"B2",  X"B4",  X"10",
  X"A0",  X"9D",  X"E0",  X"C2",  X"A0",  X"A3",  X"A4",  X"A0",
  X"80",  X"04",  X"D2",  X"83",  X"80",  X"14",  X"92",  X"7F",
  X"90",  X"80",  X"04",  X"82",  X"84",  X"C0",  X"84",  X"80",
  X"12",  X"82",  X"82",  X"83",  X"82",  X"82",  X"C8",  X"88",
  X"B4",  X"89",  X"84",  X"88",  X"02",  X"88",  X"98",  X"86",
  X"98",  X"DA",  X"9B",  X"86",  X"C6",  X"82",  X"C6",  X"84",
  X"80",  X"18",  X"87",  X"C6",  X"80",  X"A0",  X"C4",  X"C2",
  X"83",  X"C6",  X"C6",  X"A0",  X"F2",  X"E0",  X"81",  X"91",
  X"C6",  X"C6",  X"84",  X"80",  X"08",  X"82",  X"C6",  X"C6",
  X"84",  X"80",  X"18",  X"82",  X"10",  X"C4",  X"9D",  X"E0",
  X"E2",  X"80",  X"06",  X"90",  X"82",  X"A2",  X"A0",  X"C2",
  X"AC",  X"80",  X"04",  X"D2",  X"92",  X"7F",  X"AE",  X"B6",
  X"AF",  X"AE",  X"AE",  X"80",  X"1A",  X"B0",  X"82",  X"C0",
  X"82",  X"80",  X"38",  X"C0",  X"AA",  X"AB",  X"AA",  X"B2",
  X"F2",  X"B8",  X"BA",  X"B9",  X"B8",  X"B8",  X"80",  X"1A",
  X"AA",  X"23",  X"A2",  X"C2",  X"84",  X"02",  X"C4",  X"F4",
  X"A0",  X"B2",  X"E8",  X"D2",  X"40",  X"90",  X"E6",  X"D2",
  X"A4",  X"A4",  X"40",  X"91",  X"A4",  X"A7",  X"83",  X"A6",
  X"B2",  X"E4",  X"B4",  X"F2",  X"80",  X"A0",  X"18",  X"B3",
  X"F2",  X"C2",  X"83",  X"80",  X"02",  X"C2",  X"F2",  X"F4",
  X"A4",  X"A0",  X"A6",  X"E8",  X"D0",  X"92",  X"40",  X"A5",
  X"A6",  X"A6",  X"F2",  X"D0",  X"E6",  X"93",  X"40",  X"A7",
  X"A0",  X"E4",  X"B4",  X"B2",  X"80",  X"B2",  X"B2",  X"18",
  X"A7",  X"F2",  X"BA",  X"80",  X"18",  X"B6",  X"80",  X"24",
  X"EC",  X"C2",  X"80",  X"02",  X"AE",  X"EC",  X"81",  X"81",
  X"C2",  X"80",  X"32",  X"EC",  X"AC",  X"12",  X"AE",  X"EC",
  X"81",  X"81",  X"82",  X"B2",  X"10",  X"B4",  X"9D",  X"92",
  X"7F",  X"90",  X"82",  X"F2",  X"C2",  X"81",  X"91",  X"9D",
  X"E0",  X"2B",  X"A2",  X"AA",  X"A4",  X"E8",  X"92",  X"40",
  X"90",  X"93",  X"A6",  X"40",  X"90",  X"B7",  X"A6",  X"B6",
  X"83",  X"A6",  X"E6",  X"A4",  X"A2",  X"80",  X"14",  X"B7",
  X"80",  X"02",  X"01",  X"C2",  X"80",  X"36",  X"D2",  X"82",
  X"83",  X"82",  X"A0",  X"E0",  X"F6",  X"81",  X"91",  X"92",
  X"7F",  X"90",  X"D4",  X"B4",  X"92",  X"94",  X"90",  X"7F",
  X"95",  X"C4",  X"C2",  X"83",  X"C6",  X"C6",  X"F2",  X"10",
  X"B2",  X"9D",  X"82",  X"12",  X"A0",  X"B5",  X"80",  X"02",
  X"01",  X"E2",  X"80",  X"02",  X"90",  X"80",  X"12",  X"92",
  X"B5",  X"80",  X"02",  X"01",  X"D0",  X"80",  X"02",  X"92",
  X"A2",  X"80",  X"22",  X"B5",  X"92",  X"94",  X"7F",  X"90",
  X"80",  X"02",  X"B5",  X"C4",  X"C2",  X"83",  X"C6",  X"C6",
  X"F2",  X"80",  X"12",  X"B2",  X"81",  X"91",  X"94",  X"7F",
  X"90",  X"D0",  X"C0",  X"10",  X"A2",  X"82",  X"05",  X"83",
  X"84",  X"D4",  X"92",  X"90",  X"7F",  X"96",  X"10",  X"B2",
  X"7F",  X"92",  X"D0",  X"A2",  X"10",  X"C0",  X"9D",  X"92",
  X"40",  X"90",  X"A0",  X"80",  X"82",  X"04",  X"92",  X"83",
  X"80",  X"14",  X"92",  X"7F",  X"90",  X"82",  X"F8",  X"C2",
  X"80",  X"A4",  X"04",  X"A2",  X"A4",  X"D6",  X"92",  X"96",
  X"90",  X"7F",  X"94",  X"A2",  X"80",  X"34",  X"D6",  X"A4",
  X"A2",  X"A4",  X"80",  X"04",  X"B4",  X"D6",  X"92",  X"96",
  X"90",  X"7F",  X"94",  X"B4",  X"82",  X"80",  X"34",  X"D6",
  X"81",  X"91",  X"9D",  X"80",  X"12",  X"A0",  X"7F",  X"93",
  X"7F",  X"90",  X"AC",  X"C4",  X"A2",  X"80",  X"18",  X"82",
  X"A2",  X"88",  X"80",  X"1A",  X"86",  X"81",  X"91",  X"A2",
  X"86",  X"80",  X"0A",  X"89",  X"80",  X"12",  X"AE",  X"80",
  X"16",  X"A4",  X"29",  X"A8",  X"C8",  X"82",  X"80",  X"22",
  X"82",  X"EA",  X"9A",  X"9A",  X"DA",  X"80",  X"32",  X"AA",
  X"AA",  X"A4",  X"80",  X"36",  X"C8",  X"80",  X"12",  X"80",
  X"E6",  X"A6",  X"E4",  X"02",  X"A4",  X"80",  X"02",  X"84",
  X"A4",  X"80",  X"36",  X"C4",  X"A4",  X"80",  X"06",  X"92",
  X"C4",  X"C2",  X"94",  X"90",  X"C2",  X"80",  X"18",  X"C4",
  X"80",  X"82",  X"08",  X"86",  X"C4",  X"C4",  X"80",  X"86",
  X"C4",  X"C4",  X"08",  X"82",  X"C4",  X"C4",  X"80",  X"86",
  X"C4",  X"C4",  X"12",  X"82",  X"C4",  X"C4",  X"86",  X"C4",
  X"C4",  X"82",  X"C4",  X"C4",  X"B0",  X"84",  X"C8",  X"C8",
  X"C2",  X"C2",  X"10",  X"C2",  X"84",  X"B0",  X"86",  X"80",
  X"18",  X"92",  X"82",  X"82",  X"C2",  X"A4",  X"C2",  X"82",
  X"C2",  X"7F",  X"90",  X"81",  X"81",  X"82",  X"A2",  X"E2",
  X"82",  X"C2",  X"82",  X"90",  X"C4",  X"84",  X"C4",  X"7F",
  X"92",  X"30",  X"10",  X"82",  X"C6",  X"B0",  X"82",  X"C6",
  X"84",  X"10",  X"C8",  X"A4",  X"82",  X"AA",  X"80",  X"06",
  X"80",  X"C4",  X"C2",  X"94",  X"B0",  X"C2",  X"80",  X"18",
  X"C4",  X"80",  X"82",  X"08",  X"84",  X"C4",  X"C4",  X"80",
  X"84",  X"C6",  X"C6",  X"08",  X"82",  X"C4",  X"C4",  X"80",
  X"84",  X"C6",  X"C6",  X"12",  X"82",  X"C4",  X"C4",  X"84",
  X"C6",  X"C6",  X"82",  X"C6",  X"C6",  X"C6",  X"C6",  X"C2",
  X"C2",  X"82",  X"84",  X"84",  X"C4",  X"C2",  X"90",  X"C2",
  X"82",  X"A2",  X"7F",  X"E2",  X"81",  X"81",  X"92",  X"7F",
  X"90",  X"B0",  X"02",  X"84",  X"C2",  X"86",  X"86",  X"80",
  X"02",  X"94",  X"80",  X"18",  X"80",  X"84",  X"08",  X"82",
  X"C2",  X"C2",  X"80",  X"82",  X"C4",  X"C4",  X"08",  X"84",
  X"C2",  X"C2",  X"80",  X"82",  X"C4",  X"C4",  X"12",  X"84",
  X"C2",  X"C2",  X"84",  X"82",  X"C6",  X"C6",  X"C6",  X"C6",
  X"C6",  X"C6",  X"C4",  X"C4",  X"92",  X"7F",  X"90",  X"7F",
  X"90",  X"81",  X"81",  X"C2",  X"94",  X"90",  X"C2",  X"C4",
  X"80",  X"C4",  X"C2",  X"C2",  X"08",  X"C4",  X"92",  X"7F",
  X"B0",  X"84",  X"10",  X"C2",  X"EA",  X"AA",  X"9A",  X"80",
  X"06",  X"82",  X"82",  X"84",  X"84",  X"C4",  X"C2",  X"90",
  X"C2",  X"82",  X"A2",  X"7F",  X"E2",  X"81",  X"91",  X"7F",
  X"92",  X"10",  X"92",  X"10",  X"A4",  X"E4",  X"A4",  X"84",
  X"A4",  X"10",  X"B0",  X"92",  X"7F",  X"90",  X"10",  X"82",
  X"9D",  X"80",  X"02",  X"03",  X"E4",  X"80",  X"22",  X"C2",
  X"C2",  X"A0",  X"2C",  X"E4",  X"A2",  X"A3",  X"A2",  X"C2",
  X"9F",  X"A2",  X"A0",  X"3C",  X"C2",  X"E4",  X"80",  X"32",
  X"C2",  X"C2",  X"80",  X"02",  X"01",  X"9F",  X"90",  X"81",
  X"81",  X"10",  X"F0",  X"9D",  X"D2",  X"80",  X"02",  X"01",
  X"7F",  X"90",  X"7F",  X"81",  X"01",  X"9D",  X"03",  X"C2",
  X"80",  X"02",  X"01",  X"D2",  X"80",  X"22",  X"E0",  X"A2",
  X"E0",  X"80",  X"22",  X"A2",  X"92",  X"90",  X"7F",  X"E0",
  X"80",  X"12",  X"92",  X"D2",  X"A2",  X"80",  X"32",  X"E0",
  X"7F",  X"90",  X"E0",  X"80",  X"22",  X"D2",  X"A2",  X"80",
  X"22",  X"D2",  X"92",  X"90",  X"7F",  X"E0",  X"80",  X"12",
  X"92",  X"D2",  X"80",  X"22",  X"C2",  X"7F",  X"90",  X"C2",
  X"80",  X"32",  X"C2",  X"81",  X"81",  X"9F",  X"90",  X"F2",
  X"80",  X"02",  X"01",  X"7F",  X"81",  X"01",  X"82",  X"05",
  X"82",  X"09",  X"83",  X"88",  X"82",  X"82",  X"90",  X"82",
  X"91",  X"81",  X"90",  X"03",  X"82",  X"90",  X"90",  X"91",
  X"90",  X"03",  X"90",  X"81",  X"91",  X"D2",  X"03",  X"D0",
  X"82",  X"40",  X"9E",  X"01",  X"9D",  X"03",  X"D2",  X"D0",
  X"94",  X"40",  X"96",  X"80",  X"02",  X"03",  X"C4",  X"82",
  X"D0",  X"C2",  X"81",  X"91",  X"C2",  X"05",  X"82",  X"C2",
  X"81",  X"91",  X"9D",  X"C2",  X"A0",  X"80",  X"A2",  X"B6",
  X"02",  X"25",  X"D0",  X"D2",  X"94",  X"40",  X"96",  X"C2",
  X"05",  X"82",  X"F0",  X"F2",  X"C2",  X"40",  X"95",  X"01",
  X"9D",  X"03",  X"D2",  X"D0",  X"94",  X"40",  X"96",  X"80",
  X"26",  X"C2",  X"C2",  X"82",  X"C2",  X"81",  X"91",  X"05",
  X"82",  X"C2",  X"81",  X"91",  X"82",  X"80",  X"32",  X"C2",
  X"C2",  X"C4",  X"80",  X"12",  X"05",  X"07",  X"84",  X"86",
  X"88",  X"84",  X"82",  X"80",  X"22",  X"90",  X"81",  X"90",
  X"82",  X"80",  X"32",  X"90",  X"90",  X"92",  X"C2",  X"C4",
  X"80",  X"02",  X"84",  X"C2",  X"80",  X"12",  X"C6",  X"10",
  X"C2",  X"90",  X"C2",  X"92",  X"80",  X"02",  X"C6",  X"C4",
  X"80",  X"02",  X"C2",  X"86",  X"82",  X"81",  X"90",  X"C2",
  X"86",  X"82",  X"81",  X"90",  X"81",  X"01",  X"9D",  X"80",
  X"12",  X"82",  X"C2",  X"1B",  X"9A",  X"84",  X"82",  X"09",
  X"88",  X"80",  X"12",  X"82",  X"82",  X"C4",  X"86",  X"84",
  X"80",  X"32",  X"C4",  X"82",  X"C4",  X"86",  X"84",  X"80",
  X"22",  X"82",  X"10",  X"C4",  X"C4",  X"80",  X"32",  X"82",
  X"B0",  X"81",  X"81",  X"9D",  X"21",  X"90",  X"92",  X"C0",
  X"40",  X"94",  X"80",  X"02",  X"C2",  X"81",  X"91",  X"80",
  X"02",  X"01",  X"C2",  X"81",  X"91",  X"9D",  X"92",  X"40",
  X"90",  X"92",  X"7F",  X"90",  X"B0",  X"02",  X"01",  X"D4",
  X"94",  X"94",  X"80",  X"18",  X"80",  X"08",  X"82",  X"C0",
  X"C0",  X"80",  X"08",  X"82",  X"C0",  X"C0",  X"80",  X"12",
  X"82",  X"C0",  X"C0",  X"82",  X"C0",  X"C0",  X"C0",  X"81",
  X"81",  X"7F",  X"92",  X"81",  X"81",  X"9D",  X"21",  X"90",
  X"40",  X"C0",  X"80",  X"02",  X"C2",  X"81",  X"91",  X"80",
  X"02",  X"01",  X"C2",  X"81",  X"91",  X"9D",  X"80",  X"02",
  X"A0",  X"7F",  X"A4",  X"C2",  X"80",  X"02",  X"01",  X"23",
  X"D0",  X"80",  X"22",  X"C2",  X"C2",  X"80",  X"02",  X"01",
  X"C2",  X"83",  X"80",  X"02",  X"83",  X"80",  X"12",  X"A0",
  X"C2",  X"80",  X"22",  X"C2",  X"9F",  X"D0",  X"80",  X"26",
  X"A0",  X"C2",  X"80",  X"32",  X"D2",  X"D2",  X"80",  X"02",
  X"82",  X"80",  X"22",  X"C0",  X"7F",  X"D0",  X"C0",  X"D2",
  X"80",  X"22",  X"C0",  X"7F",  X"D0",  X"C0",  X"C0",  X"40",
  X"90",  X"40",  X"90",  X"7F",  X"01",  X"81",  X"91",  X"40",
  X"90",  X"10",  X"23",  X"40",  X"90",  X"7F",  X"A0",  X"81",
  X"91",  X"7F",  X"01",  X"C2",  X"83",  X"80",  X"12",  X"83",
  X"30",  X"7F",  X"90",  X"10",  X"D2",  X"7F",  X"90",  X"10",
  X"A0",  X"92",  X"03",  X"D0",  X"82",  X"7F",  X"9E",  X"01",
  X"9D",  X"21",  X"90",  X"92",  X"40",  X"C0",  X"80",  X"02",
  X"C2",  X"81",  X"91",  X"80",  X"02",  X"01",  X"C2",  X"81",
  X"91",  X"9D",  X"21",  X"90",  X"92",  X"C0",  X"40",  X"94",
  X"80",  X"02",  X"C2",  X"81",  X"91",  X"80",  X"02",  X"01",
  X"C2",  X"81",  X"91",  X"9D",  X"21",  X"90",  X"92",  X"C0",
  X"40",  X"94",  X"80",  X"02",  X"C2",  X"81",  X"91",  X"80",
  X"02",  X"01",  X"C2",  X"81",  X"91",  X"98",  X"81",  X"9A",
  X"02",  X"98",  X"99",  X"99",  X"99",  X"99",  X"99",  X"99",
  X"99",  X"99",  X"99",  X"99",  X"99",  X"99",  X"99",  X"99",
  X"99",  X"99",  X"99",  X"99",  X"99",  X"99",  X"99",  X"99",
  X"99",  X"99",  X"99",  X"99",  X"99",  X"99",  X"99",  X"99",
  X"99",  X"99",  X"99",  X"81",  X"91",  X"99",  X"99",  X"99",
  X"99",  X"99",  X"99",  X"99",  X"99",  X"99",  X"99",  X"99",
  X"99",  X"99",  X"9B",  X"99",  X"9B",  X"81",  X"90",  X"10",
  X"86",  X"80",  X"16",  X"86",  X"80",  X"16",  X"80",  X"16",
  X"92",  X"90",  X"9A",  X"12",  X"96",  X"91",  X"81",  X"90",
  X"80",  X"0A",  X"94",  X"03",  X"80",  X"0A",  X"98",  X"80",
  X"1A",  X"84",  X"9B",  X"10",  X"98",  X"9A",  X"1A",  X"84",
  X"83",  X"9B",  X"9A",  X"10",  X"84",  X"80",  X"0A",  X"01",
  X"02",  X"01",  X"84",  X"06",  X"01",  X"96",  X"94",  X"10",
  X"01",  X"95",  X"06",  X"9B",  X"96",  X"10",  X"94",  X"96",
  X"94",  X"84",  X"16",  X"80",  X"30",  X"9B",  X"80",  X"08",
  X"98",  X"02",  X"98",  X"80",  X"95",  X"06",  X"9B",  X"96",
  X"06",  X"9B",  X"96",  X"06",  X"9B",  X"96",  X"06",  X"9B",
  X"96",  X"10",  X"94",  X"96",  X"10",  X"94",  X"96",  X"06",
  X"9B",  X"96",  X"10",  X"94",  X"96",  X"10",  X"94",  X"96",
  X"06",  X"9B",  X"96",  X"06",  X"9B",  X"96",  X"10",  X"94",
  X"96",  X"10",  X"94",  X"96",  X"06",  X"9B",  X"96",  X"10",
  X"94",  X"96",  X"10",  X"94",  X"96",  X"06",  X"9B",  X"96",
  X"06",  X"9B",  X"96",  X"06",  X"9B",  X"96",  X"10",  X"94",
  X"96",  X"10",  X"94",  X"96",  X"06",  X"9B",  X"96",  X"10",
  X"94",  X"96",  X"10",  X"94",  X"96",  X"06",  X"9B",  X"96",
  X"06",  X"9B",  X"96",  X"10",  X"94",  X"96",  X"10",  X"94",
  X"96",  X"06",  X"9B",  X"96",  X"10",  X"94",  X"96",  X"10",
  X"94",  X"98",  X"16",  X"80",  X"26",  X"94",  X"80",  X"26",
  X"94",  X"81",  X"90",  X"10",  X"86",  X"80",  X"16",  X"86",
  X"80",  X"16",  X"80",  X"16",  X"92",  X"90",  X"9A",  X"12",
  X"96",  X"91",  X"81",  X"90",  X"80",  X"0A",  X"94",  X"03",
  X"80",  X"0A",  X"98",  X"80",  X"1A",  X"84",  X"9B",  X"10",
  X"98",  X"9A",  X"1A",  X"84",  X"83",  X"9B",  X"9A",  X"10",
  X"84",  X"80",  X"0A",  X"01",  X"02",  X"01",  X"84",  X"06",
  X"01",  X"96",  X"94",  X"10",  X"01",  X"95",  X"06",  X"9B",
  X"96",  X"10",  X"94",  X"96",  X"94",  X"84",  X"16",  X"80",
  X"30",  X"9B",  X"80",  X"08",  X"98",  X"02",  X"98",  X"80",
  X"95",  X"06",  X"9B",  X"96",  X"06",  X"9B",  X"96",  X"06",
  X"9B",  X"96",  X"06",  X"9B",  X"96",  X"10",  X"94",  X"96",
  X"10",  X"94",  X"96",  X"06",  X"9B",  X"96",  X"10",  X"94",
  X"96",  X"10",  X"94",  X"96",  X"06",  X"9B",  X"96",  X"06",
  X"9B",  X"96",  X"10",  X"94",  X"96",  X"10",  X"94",  X"96",
  X"06",  X"9B",  X"96",  X"10",  X"94",  X"96",  X"10",  X"94",
  X"96",  X"06",  X"9B",  X"96",  X"06",  X"9B",  X"96",  X"06",
  X"9B",  X"96",  X"10",  X"94",  X"96",  X"10",  X"94",  X"96",
  X"06",  X"9B",  X"96",  X"10",  X"94",  X"96",  X"10",  X"94",
  X"96",  X"06",  X"9B",  X"96",  X"06",  X"9B",  X"96",  X"10",
  X"94",  X"96",  X"10",  X"94",  X"96",  X"06",  X"9B",  X"96",
  X"10",  X"94",  X"96",  X"10",  X"94",  X"98",  X"16",  X"80",
  X"26",  X"96",  X"80",  X"26",  X"96",  X"81",  X"90",  X"81",
  X"90",  X"03",  X"90",  X"C2",  X"81",  X"C0",  X"81",  X"90",
  X"9D",  X"40",  X"B0",  X"82",  X"C2",  X"81",  X"81",  X"9D",
  X"80",  X"14",  X"B0",  X"30",  X"02",  X"01",  X"B0",  X"80",
  X"04",  X"01",  X"40",  X"01",  X"D0",  X"91",  X"91",  X"80",
  X"12",  X"80",  X"81",  X"91",  X"81",  X"81",  X"05",  X"C2",
  X"80",  X"22",  X"03",  X"90",  X"D0",  X"81",  X"90",  X"82",
  X"90",  X"C2",  X"D0",  X"81",  X"90",  X"9D",  X"80",  X"04",
  X"A0",  X"10",  X"D0",  X"40",  X"91",  X"A0",  X"80",  X"04",
  X"01",  X"D0",  X"91",  X"83",  X"80",  X"12",  X"01",  X"40",
  X"90",  X"D0",  X"91",  X"40",  X"91",  X"A0",  X"80",  X"34",
  X"D0",  X"81",  X"91",  X"03",  X"C2",  X"86",  X"C4",  X"80",
  X"02",  X"84",  X"C4",  X"80",  X"02",  X"01",  X"81",  X"01",
  X"C4",  X"80",  X"02",  X"84",  X"C4",  X"81",  X"01",  X"03",
  X"C6",  X"80",  X"84",  X"02",  X"90",  X"C2",  X"80",  X"02",
  X"01",  X"D0",  X"81",  X"01",  X"A7",  X"AE",  X"83",  X"29",
  X"E8",  X"A9",  X"82",  X"81",  X"81",  X"01",  X"01",  X"01",
  X"E0",  X"E4",  X"E8",  X"EC",  X"F0",  X"F4",  X"F8",  X"FC",
  X"81",  X"82",  X"81",  X"81",  X"01",  X"01",  X"01",  X"A7",
  X"A9",  X"2B",  X"EA",  X"AB",  X"AA",  X"81",  X"01",  X"01",
  X"01",  X"81",  X"81",  X"E0",  X"E4",  X"E8",  X"EC",  X"F0",
  X"F4",  X"F8",  X"FC",  X"81",  X"81",  X"81",  X"81",  X"A7",
  X"29",  X"AD",  X"01",  X"27",  X"A6",  X"E0",  X"81",  X"01",
  X"01",  X"01",  X"9D",  X"9D",  X"9D",  X"9D",  X"9D",  X"9D",
  X"9D",  X"81",  X"81",  X"81",  X"81",  X"81",  X"81",  X"81",
  X"27",  X"A6",  X"C0",  X"E2",  X"A4",  X"E2",  X"E4",  X"10",
  X"AC",  X"29",  X"A8",  X"C2",  X"C8",  X"E0",  X"E2",  X"E4",
  X"E8",  X"81",  X"83",  X"82",  X"81",  X"01",  X"01",  X"01",
  X"09",  X"C8",  X"81",  X"88",  X"80",  X"02",  X"01",  X"01",
  X"80",  X"12",  X"01",  X"09",  X"C8",  X"81",  X"80",  X"02",
  X"01",  X"01",  X"88",  X"80",  X"12",  X"01",  X"81",  X"29",
  X"A8",  X"C8",  X"C2",  X"E0",  X"E2",  X"E4",  X"C0",  X"81",
  X"01",  X"01",  X"01",  X"81",  X"81",  X"A0",  X"81",  X"01",
  X"01",  X"01",  X"81",  X"81",  X"80",  X"12",  X"A8",  X"81",
  X"B0",  X"30",  X"80",  X"12",  X"A8",  X"AA",  X"A8",  X"81",
  X"30",  X"80",  X"12",  X"A9",  X"A8",  X"81",  X"01",  X"01",
  X"01",  X"30",  X"80",  X"12",  X"A9",  X"A8",  X"81",  X"01",
  X"01",  X"01",  X"30",  X"80",  X"12",  X"01",  X"30",  X"91",
  X"81",  X"81",  X"92",  X"81",  X"91",  X"92",  X"81",  X"91",
  X"92",  X"81",  X"91",  X"27",  X"A0",  X"A6",  X"81",  X"01",
  X"01",  X"01",  X"A7",  X"29",  X"A6",  X"12",  X"01",  X"91",
  X"29",  X"A8",  X"E8",  X"2B",  X"AA",  X"EA",  X"80",  X"02",
  X"01",  X"80",  X"02",  X"01",  X"C1",  X"C5",  X"C9",  X"CD",
  X"D1",  X"D5",  X"D9",  X"DD",  X"E1",  X"E5",  X"E9",  X"ED",
  X"F1",  X"F5",  X"F9",  X"FD",  X"C1",  X"2D",  X"AC",  X"E8",
  X"80",  X"02",  X"01",  X"C1",  X"C5",  X"C9",  X"CD",  X"D1",
  X"D5",  X"D9",  X"DD",  X"E1",  X"E5",  X"E9",  X"ED",  X"F1",
  X"F5",  X"F9",  X"FD",  X"C1",  X"81",  X"01",  X"01",  X"01",
  X"81",  X"81",  X"81",  X"01",  X"81",  X"01",  X"81",  X"01",
  X"AE",  X"A7",  X"2D",  X"AC",  X"29",  X"81",  X"01",  X"11",
  X"90",  X"D2",  X"92",  X"D2",  X"93",  X"90",  X"92",  X"11",
  X"90",  X"D0",  X"80",  X"22",  X"92",  X"81",  X"01",  X"01",
  X"01",  X"90",  X"40",  X"92",  X"92",  X"81",  X"01",  X"01",
  X"01",  X"11",  X"90",  X"D2",  X"92",  X"D2",  X"10",  X"AC",
  X"9D",  X"1B",  X"89",  X"9A",  X"80",  X"82",  X"14",  X"C6",
  X"B3",  X"19",  X"80",  X"98",  X"02",  X"84",  X"80",  X"12",
  X"82",  X"10",  X"C2",  X"22",  X"C2",  X"C2",  X"80",  X"12",
  X"80",  X"C4",  X"F0",  X"C6",  X"82",  X"81",  X"91",  X"F0",
  X"81",  X"91",  X"91",  X"03",  X"82",  X"C4",  X"C4",  X"81",
  X"D2",  X"9D",  X"05",  X"82",  X"C2",  X"80",  X"22",  X"C4",
  X"80",  X"22",  X"B0",  X"A3",  X"03",  X"82",  X"E0",  X"80",
  X"02",  X"29",  X"2D",  X"2B",  X"27",  X"A8",  X"AC",  X"AA",
  X"10",  X"A6",  X"A4",  X"84",  X"C4",  X"C4",  X"80",  X"22",
  X"D2",  X"9F",  X"01",  X"C2",  X"D2",  X"90",  X"9F",  X"94",
  X"C2",  X"80",  X"22",  X"C2",  X"9F",  X"01",  X"C2",  X"82",
  X"C2",  X"E0",  X"80",  X"02",  X"01",  X"C2",  X"80",  X"22",
  X"E0",  X"C4",  X"80",  X"12",  X"C4",  X"80",  X"02",  X"A4",
  X"E0",  X"80",  X"32",  X"C2",  X"81",  X"81",  X"F0",  X"10",
  X"B0",  X"8C",  X"A7",  X"8B",  X"8A",  X"80",  X"02",  X"0B",
  X"8A",  X"09",  X"88",  X"C8",  X"0B",  X"8A",  X"09",  X"88",
  X"C8",  X"10",  X"90",  X"92",  X"40",  X"01",  X"80",  X"02",
  X"01",  X"C2",  X"11",  X"82",  X"11",  X"84",  X"90",  X"92",
  X"94",  X"40",  X"01",  X"80",  X"02",  X"01",  X"40",  X"92",
  X"0B",  X"8A",  X"D2",  X"90",  X"92",  X"94",  X"40",  X"01",
  X"80",  X"02",  X"01",  X"40",  X"92",  X"92",  X"0B",  X"8A",
  X"D2",  X"90",  X"92",  X"94",  X"40",  X"01",  X"80",  X"02",
  X"01",  X"40",  X"92",  X"0B",  X"8A",  X"D2",  X"D4",  X"95",
  X"94",  X"D4",  X"9E",  X"81",  X"01",  X"03",  X"82",  X"82",
  X"91",  X"81",  X"01",  X"9D",  X"03",  X"C2",  X"84",  X"80",
  X"02",  X"B0",  X"90",  X"9F",  X"92",  X"B0",  X"81",  X"81",
  X"9D",  X"03",  X"C2",  X"80",  X"02",  X"84",  X"9F",  X"90",
  X"84",  X"81",  X"91",  X"9D",  X"03",  X"C2",  X"80",  X"02",
  X"84",  X"9F",  X"90",  X"84",  X"81",  X"91",  X"9D",  X"03",
  X"C2",  X"80",  X"02",  X"84",  X"9F",  X"90",  X"84",  X"81",
  X"91",  X"9D",  X"03",  X"C2",  X"80",  X"02",  X"84",  X"9F",
  X"90",  X"84",  X"81",  X"91",  X"9D",  X"03",  X"C2",  X"80",
  X"02",  X"84",  X"9F",  X"90",  X"84",  X"81",  X"91",  X"9D",
  X"03",  X"C2",  X"80",  X"02",  X"84",  X"9F",  X"90",  X"84",
  X"81",  X"91",  X"9D",  X"03",  X"C2",  X"84",  X"80",  X"02",
  X"B0",  X"90",  X"9F",  X"92",  X"B0",  X"81",  X"81",  X"01",
  X"03",  X"82",  X"9F",  X"01",  X"03",  X"82",  X"81",  X"03",
  X"82",  X"9F",  X"01",  X"03",  X"82",  X"9F",  X"01",  X"8B",
  X"8B",  X"8A",  X"80",  X"12",  X"01",  X"8B",  X"8B",  X"80",
  X"12",  X"01",  X"7F",  X"01",  X"7F",  X"01",  X"9C",  X"7F",
  X"01",  X"82",  X"91",  X"01",  X"29",  X"A6",  X"32",  X"A0",
  X"91",  X"81",  X"01",  X"01",  X"01",  X"81",  X"81",  X"81",
  X"01",  X"81",  X"01",  X"A7",  X"8B",  X"8A",  X"80",  X"12",
  X"01",  X"21",  X"A0",  X"A2",  X"E2",  X"8B",  X"10",  X"21",
  X"A0",  X"A2",  X"E2",  X"21",  X"E6",  X"8B",  X"8A",  X"27",
  X"A6",  X"CA",  X"8A",  X"27",  X"A6",  X"CA",  X"27",  X"A6",
  X"8A",  X"CA",  X"81",  X"01",  X"81",  X"01",  X"91",  X"01",
  X"01",  X"01",  X"81",  X"81",  X"83",  X"83",  X"82",  X"80",
  X"12",  X"01",  X"83",  X"05",  X"82",  X"A3",  X"88",  X"09",
  X"81",  X"01",  X"9D",  X"21",  X"23",  X"A0",  X"A2",  X"80",
  X"1A",  X"01",  X"D0",  X"80",  X"02",  X"A0",  X"9F",  X"01",
  X"80",  X"2A",  X"D0",  X"81",  X"81",  X"AA",  X"E0",  X"E2",
  X"E4",  X"C2",  X"C4",  X"C8",  X"CC",  X"85",  X"C4",  X"F0",
  X"F4",  X"F8",  X"FC",  X"05",  X"C6",  X"C6",  X"86",  X"C6",
  X"A8",  X"A9",  X"80",  X"02",  X"01",  X"85",  X"07",  X"C6",
  X"A7",  X"84",  X"84",  X"81",  X"81",  X"E0",  X"E4",  X"E8",
  X"EC",  X"F0",  X"F4",  X"F8",  X"FC",  X"81",  X"81",  X"9C",
  X"05",  X"84",  X"C4",  X"80",  X"02",  X"01",  X"9F",  X"92",
  X"C4",  X"07",  X"C4",  X"81",  X"82",  X"83",  X"05",  X"C4",
  X"85",  X"82",  X"85",  X"80",  X"02",  X"83",  X"07",  X"C6",
  X"85",  X"82",  X"82",  X"81",  X"C2",  X"81",  X"F0",  X"F4",
  X"F8",  X"FC",  X"C2",  X"C4",  X"C8",  X"CC",  X"E0",  X"E2",
  X"E4",  X"81",  X"E0",  X"E4",  X"E8",  X"EC",  X"F0",  X"F4",
  X"F8",  X"FC",  X"10",  X"81",  X"C2",  X"81",  X"F0",  X"F4",
  X"F8",  X"FC",  X"C2",  X"C4",  X"C8",  X"CC",  X"E0",  X"E2",
  X"E4",  X"81",  X"01",  X"01",  X"01",  X"81",  X"81",  X"AA",
  X"E0",  X"29",  X"A0",  X"C2",  X"C4",  X"C8",  X"CC",  X"85",
  X"C4",  X"05",  X"C6",  X"C6",  X"86",  X"C6",  X"C0",  X"A8",
  X"A9",  X"80",  X"02",  X"01",  X"85",  X"07",  X"C6",  X"A7",
  X"84",  X"84",  X"81",  X"81",  X"E0",  X"E4",  X"E8",  X"EC",
  X"F0",  X"F4",  X"F8",  X"FC",  X"81",  X"81",  X"9C",  X"05",
  X"84",  X"C4",  X"80",  X"02",  X"01",  X"9F",  X"92",  X"C4",
  X"07",  X"C4",  X"07",  X"C6",  X"80",  X"12",  X"01",  X"C4",
  X"07",  X"84",  X"A0",  X"A0",  X"30",  X"84",  X"80",  X"12",
  X"07",  X"C0",  X"81",  X"82",  X"83",  X"05",  X"C4",  X"85",
  X"82",  X"85",  X"80",  X"02",  X"83",  X"07",  X"C6",  X"85",
  X"82",  X"82",  X"81",  X"C2",  X"81",  X"C2",  X"C4",  X"C8",
  X"CC",  X"81",  X"E0",  X"E4",  X"E8",  X"EC",  X"F0",  X"F4",
  X"F8",  X"FC",  X"10",  X"81",  X"C2",  X"81",  X"C2",  X"C4",
  X"C8",  X"CC",  X"81",  X"01",  X"01",  X"01",  X"81",  X"81",
  X"82",  X"9A",  X"96",  X"91",  X"98",  X"D4",  X"91",  X"80",
  X"32",  X"96",  X"91",  X"90",  X"80",  X"02",  X"94",  X"96",
  X"80",  X"28",  X"91",  X"94",  X"81",  X"90",  X"82",  X"98",
  X"91",  X"9A",  X"D6",  X"91",  X"80",  X"32",  X"98",  X"91",
  X"90",  X"80",  X"02",  X"96",  X"98",  X"80",  X"28",  X"91",
  X"96",  X"81",  X"90",  X"D4",  X"17",  X"92",  X"90",  X"91",
  X"92",  X"11",  X"90",  X"94",  X"95",  X"94",  X"92",  X"81",
  X"90",  X"03",  X"81",  X"D0",  X"9D",  X"21",  X"A0",  X"C2",
  X"80",  X"02",  X"A0",  X"9F",  X"A0",  X"C2",  X"80",  X"12",
  X"01",  X"81",  X"81",  X"9D",  X"81",  X"81",  X"00",  X"00",
  X"00",  X"00",  X"01",  X"04",  X"1B",  X"00",  X"00",  X"FF",
  X"00",  X"00",  X"00",  X"00",  X"01",  X"00",  X"06",  X"C5",
  X"0E",  X"00",  X"00",  X"FF",  X"00",  X"00",  X"2D",  X"1F",
  X"00",  X"00",  X"FF",  X"00",  X"00",  X"2D",  X"1F",  X"00",
  X"00",  X"FF",  X"00",  X"00",  X"2D",  X"1F",  X"00",  X"00",
  X"FF",  X"00",  X"00",  X"2D",  X"1F",  X"00",  X"00",  X"FF",
  X"00",  X"00",  X"2D",  X"1F",  X"00",  X"00",  X"FF",  X"00",
  X"00",  X"2D",  X"1F",  X"00",  X"00",  X"FF",  X"00",  X"00",
  X"2D",  X"1F",  X"00",  X"00",  X"FF",  X"00",  X"00",  X"2D",
  X"1F",  X"00",  X"00",  X"FF",  X"00",  X"00",  X"2D",  X"1F",
  X"00",  X"00",  X"FF",  X"00",  X"00",  X"2D",  X"1F",  X"00",
  X"00",  X"FF",  X"00",  X"00",  X"2D",  X"1F",  X"00",  X"00",
  X"FF",  X"00",  X"00",  X"00",  X"00",  X"FF",  X"00",  X"00",
  X"2D",  X"1F",  X"00",  X"00",  X"FF",  X"00",  X"00",  X"2D",
  X"1F",  X"00",  X"00",  X"FF",  X"00",  X"00",  X"2D",  X"1F",
  X"00",  X"00",  X"FF",  X"00",  X"00",  X"00",  X"00",  X"FF",
  X"00",  X"00",  X"00",  X"00",  X"FF",  X"00",  X"00",  X"2D",
  X"1F",  X"00",  X"00",  X"FF",  X"00",  X"00",  X"00",  X"00",
  X"FF",  X"00",  X"00",  X"00",  X"00",  X"FF",  X"00",  X"00",
  X"2D",  X"1F",  X"00",  X"00",  X"FF",  X"00",  X"00",  X"2D",
  X"1F",  X"00",  X"00",  X"FF",  X"00",  X"00",  X"2D",  X"00",
  X"00",  X"FF",  X"00",  X"00",  X"00",  X"00",  X"FF",  X"00",
  X"00",  X"2D",  X"1F",  X"00",  X"00",  X"FF",  X"00",  X"00",
  X"00",  X"00",  X"FF",  X"00",  X"00",  X"2D",  X"1F",  X"00",
  X"00",  X"FF",  X"00",  X"00",  X"00",  X"00",  X"FF",  X"00",
  X"00",  X"2D",  X"1F",  X"00",  X"00",  X"FF",  X"00",  X"00",
  X"2D",  X"1F",  X"00",  X"00",  X"FF",  X"00",  X"00",  X"2D",
  X"1F",  X"00",  X"00",  X"FF",  X"00",  X"00",  X"2D",  X"1F",
  X"00",  X"00",  X"FF",  X"00",  X"00",  X"2D",  X"1F",  X"00",
  X"00",  X"FF",  X"00",  X"00",  X"00",  X"00",  X"FF",  X"00",
  X"00",  X"00",  X"00",  X"FF",  X"00",  X"00",  X"2D",  X"1F",
  X"00",  X"00",  X"FF",  X"00",  X"00",  X"00",  X"00",  X"FF",
  X"00",  X"00",  X"2D",  X"1F",  X"00",  X"00",  X"FF",  X"00",
  X"00",  X"2D",  X"1F",  X"00",  X"00",  X"FF",  X"00",  X"00",
  X"00",  X"00",  X"FF",  X"00",  X"00",  X"2D",  X"00",  X"00",
  X"FF",  X"00",  X"00",  X"2D",  X"1F",  X"00",  X"00",  X"FF",
  X"00",  X"00",  X"2D",  X"1F",  X"00",  X"00",  X"FF",  X"00",
  X"00",  X"2D",  X"1F",  X"00",  X"00",  X"FF",  X"00",  X"00",
  X"2D",  X"00",  X"00",  X"FF",  X"00",  X"00",  X"2D",  X"00",
  X"00",  X"FF",  X"00",  X"00",  X"2D",  X"1F",  X"00",  X"00",
  X"FF",  X"00",  X"00",  X"2D",  X"1F",  X"00",  X"00",  X"FF",
  X"00",  X"00",  X"2D",  X"00",  X"00",  X"FF",  X"00",  X"00",
  X"2D",  X"00",  X"00",  X"FF",  X"00",  X"00",  X"00",  X"00",
  X"FF",  X"00",  X"00",  X"00",  X"00",  X"FF",  X"00",  X"00",
  X"00",  X"00",  X"FF",  X"00",  X"00",  X"2D",  X"1F",  X"00",
  X"00",  X"FF",  X"00",  X"00",  X"00",  X"00",  X"FF",  X"00",
  X"00",  X"2D",  X"1F",  X"00",  X"00",  X"FF",  X"00",  X"00",
  X"2D",  X"1F",  X"00",  X"00",  X"FF",  X"00",  X"00",  X"2D",
  X"1F",  X"00",  X"00",  X"FF",  X"00",  X"00",  X"2D",  X"1F",
  X"00",  X"00",  X"FF",  X"00",  X"00",  X"2D",  X"1F",  X"00",
  X"00",  X"FF",  X"00",  X"00",  X"00",  X"00",  X"FF",  X"00",
  X"00",  X"00",  X"00",  X"FF",  X"00",  X"00",  X"00",  X"00",
  X"FF",  X"00",  X"00",  X"2D",  X"1F",  X"00",  X"00",  X"FF",
  X"00",  X"00",  X"00",  X"00",  X"FF",  X"00",  X"00",  X"2D",
  X"1F",  X"00",  X"00",  X"FF",  X"00",  X"00",  X"2D",  X"1F",
  X"00",  X"00",  X"FF",  X"00",  X"00",  X"00",  X"00",  X"FF",
  X"00",  X"00",  X"2D",  X"1F",  X"00",  X"00",  X"FF",  X"00",
  X"00",  X"2D",  X"1F",  X"00",  X"00",  X"FF",  X"00",  X"00",
  X"2D",  X"1F",  X"00",  X"00",  X"FF",  X"00",  X"00",  X"2D",
  X"1F",  X"00",  X"00",  X"FF",  X"00",  X"00",  X"2D",  X"1F",
  X"00",  X"00",  X"FF",  X"00",  X"00",  X"2D",  X"1F",  X"00",
  X"00",  X"FF",  X"00",  X"00",  X"2D",  X"1F",  X"00",  X"00",
  X"FF",  X"00",  X"00",  X"2D",  X"1F",  X"00",  X"00",  X"FF",
  X"00",  X"00",  X"2D",  X"1F",  X"00",  X"00",  X"FF",  X"00",
  X"00",  X"2D",  X"1F",  X"00",  X"00",  X"FF",  X"00",  X"00",
  X"2D",  X"1F",  X"00",  X"00",  X"FF",  X"00",  X"00",  X"2D",
  X"1F",  X"00",  X"00",  X"FF",  X"00",  X"00",  X"2D",  X"1F",
  X"00",  X"00",  X"FF",  X"00",  X"00",  X"00",  X"00",  X"FF",
  X"00",  X"00",  X"00",  X"00",  X"FF",  X"00",  X"00",  X"00",
  X"00",  X"FF",  X"00",  X"00",  X"2D",  X"1F",  X"00",  X"00",
  X"FF",  X"00",  X"00",  X"2D",  X"1F",  X"00",  X"00",  X"FF",
  X"00",  X"00",  X"2D",  X"1F",  X"00",  X"00",  X"FF",  X"00",
  X"00",  X"00",  X"00",  X"FF",  X"00",  X"00",  X"2D",  X"1F",
  X"00",  X"00",  X"FF",  X"00",  X"00",  X"2D",  X"1F",  X"00",
  X"00",  X"FF",  X"00",  X"00",  X"2D",  X"1F",  X"00",  X"00",
  X"FF",  X"00",  X"00",  X"2D",  X"1F",  X"00",  X"00",  X"FF",
  X"00",  X"00",  X"2D",  X"1F",  X"00",  X"00",  X"FF",  X"00",
  X"00",  X"00",  X"00",  X"FF",  X"00",  X"00",  X"2D",  X"1F",
  X"00",  X"00",  X"FF",  X"00",  X"00",  X"2D",  X"1F",  X"00",
  X"00",  X"FF",  X"00",  X"00",  X"2D",  X"1F",  X"00",  X"00",
  X"FF",  X"00",  X"00",  X"00",  X"00",  X"FF",  X"00",  X"00",
  X"00",  X"00",  X"FF",  X"00",  X"00",  X"00",  X"00",  X"FF",
  X"00",  X"00",  X"2D",  X"00",  X"00",  X"FF",  X"00",  X"00",
  X"2D",  X"1F",  X"00",  X"00",  X"FF",  X"00",  X"00",  X"00",
  X"00",  X"FF",  X"00",  X"00",  X"2D",  X"1F",  X"00",  X"00",
  X"FF",  X"00",  X"00",  X"00",  X"00",  X"FF",  X"00",  X"00",
  X"00",  X"00",  X"FF",  X"00",  X"00",  X"2D",  X"1F",  X"00",
  X"00",  X"FF",  X"00",  X"00",  X"00",  X"00",  X"FF",  X"00",
  X"00",  X"2D",  X"1F",  X"00",  X"00",  X"FF",  X"00",  X"00",
  X"00",  X"00",  X"FF",  X"00",  X"00",  X"2D",  X"1F",  X"00",
  X"00",  X"FF",  X"00",  X"00",  X"2D",  X"1F",  X"00",  X"00",
  X"FF",  X"00",  X"00",  X"2D",  X"1F",  X"00",  X"00",  X"FF",
  X"00",  X"00",  X"2D",  X"1F",  X"00",  X"00",  X"FF",  X"00",
  X"00",  X"2D",  X"1F",  X"00",  X"00",  X"FF",  X"00",  X"00",
  X"2D",  X"1F",  X"00",  X"00",  X"FF",  X"00",  X"00",  X"2D",
  X"1F",  X"00",  X"00",  X"FF",  X"00",  X"00",  X"2D",  X"1F",
  X"00",  X"00",  X"FF",  X"00",  X"00",  X"2D",  X"1F",  X"00",
  X"00",  X"FF",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"FF",  X"00",  X"00",  X"00",  X"FF",  X"00",  X"00",
  X"80",  X"80",  X"80",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"80",  X"80",  X"80",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"25",  X"25",  X"49",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"80",  X"80",  X"80",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"80",  X"80",  X"80",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"40",  X"51",  X"80",  X"80",
  X"80",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"40",  X"00",  X"43",  X"00",  X"30",  X"34",
  X"38",  X"43",  X"00",  X"00",  X"49",  X"00",  X"30",  X"34",
  X"38",  X"63",  X"00",  X"00",  X"4E",  X"00",  X"30",  X"00",
  X"2E",  X"00",  X"28",  X"6C",  X"00",  X"00",  X"30",  X"30",
  X"30",  X"30",  X"20",  X"20",  X"20",  X"20",  X"43",  X"46",
  X"43",  X"49",  X"43",  X"43",  X"43",  X"53",  X"49",  X"6E",
  X"00",  X"00",  X"41",  X"00",  X"3F",  X"00",  X"3F",  X"63",
  X"3F",  X"8B",  X"3F",  X"50",  X"3F",  X"00",  X"40",  X"00",
  X"40",  X"00",  X"40",  X"00",  X"3F",  X"00",  X"49",  X"38",
  X"2D",  X"00",  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",
  X"40",  X"40",  X"40",  X"40",  X"7F",  X"7F",  X"40",  X"00",
  X"3F",  X"00",  X"40",  X"00",  X"40",  X"00",  X"40",  X"00",
  X"40",  X"00",  X"40",  X"00",  X"41",  X"00",  X"41",  X"00",
  X"41",  X"00",  X"41",  X"00",  X"42",  X"20",  X"42",  X"E8",
  X"42",  X"A2",  X"42",  X"E5",  X"42",  X"1E",  X"43",  X"26",
  X"43",  X"37",  X"43",  X"85",  X"43",  X"67",  X"43",  X"60",
  X"44",  X"78",  X"44",  X"D6",  X"44",  X"06",  X"44",  X"C7",
  X"44",  X"79",  X"43",  X"37",  X"46",  X"B5",  X"4D",  X"E9",
  X"5A",  X"F9",  X"75",  X"7F",  X"3C",  X"97",  X"39",  X"D5",
  X"32",  X"44",  X"25",  X"CF",  X"0A",  X"64",  X"00",  X"00",
  X"00",  X"00",  X"9D",  X"7F",  X"01",  X"7F",  X"01",  X"81",
  X"81",  X"9D",  X"7F",  X"01",  X"81",  X"81",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"40",  X"00",  X"00",  X"40",
  X"40",  X"40",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"40",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"33",  X"12",  X"DE",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"40",  X"40",  X"40",  X"40",
  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",
  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",
  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",
  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",
  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",
  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",
  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",
  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",
  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",
  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",
  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",
  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",
  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",
  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",
  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",
  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",
  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",
  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",
  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",
  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",
  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",
  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",
  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",
  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",
  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",
  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",
  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",
  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",
  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",
  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",
  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",  X"40",
  X"40",  X"40",  X"40",  X"40",  X"00",  X"FF",  X"00",  X"40",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"40",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"43",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"40",  X"40",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"80",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"FF",  X"80",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",  X"00",
  others => X"00" );



end;
