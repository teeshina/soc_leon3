----------------------------------------------------------------------------
--  INFORMATION:  http://www.GNSS-sensor.com
--  PROPERTY:     GNSS Sensor Ltd
--  E-MAIL:       alex.kosin@gnss-sensor.com
--  DESCRIPTION:  This file contains copy of firmware image
------------------------------------------------------------------------------
--  WARNING:      
------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
library grlib;
use grlib.amba.all;
use grlib.stdlib.all;
--use grlib.devices.all;

entity FwRomImage is
  generic (
    hindex  : integer := 0;
    haddr   : integer := 0;
    hmask   : integer := 16#fff#);
  port (
    rst     : in  std_ulogic;
    clk     : in  std_ulogic;
    ahbsi   : in  ahb_slv_in_type;
    ahbso   : out ahb_slv_out_type
  );
end;

architecture rtl of FwRomImage is

constant VENDOR_GNSSSENSOR     : integer := 16#F1#; -- TODO: move to devices.vhd
constant GNSSSENSOR_ROM_IMAGE  : integer := 16#07B#;
constant REVISION              : integer := 1;

constant hconfig : ahb_config_type := (
  0 => ahb_device_reg ( VENDOR_GNSSSENSOR, GNSSSENSOR_ROM_IMAGE, 0, REVISION, 0),
  4 => ahb_membar(haddr, '1', '1', hmask), others => zero32);

signal romdata : std_logic_vector(31 downto 0);
signal addr : std_logic_vector(15 downto 0);
signal hsel, hready : std_ulogic;

begin

  ahbso.hresp   <= "00";
  ahbso.hsplit  <= (others => '0');
  ahbso.hirq    <= (others => '0');
  ahbso.hcache  <= '1';
  ahbso.hconfig <= hconfig;
  ahbso.hindex  <= hindex;
  
  reg : process (clk) begin
    if rising_edge(clk) then addr <= ahbsi.haddr(17 downto 2); end if;
  end process;
  
  ahbso.hrdata  <= romdata;
  ahbso.hready  <= '1';
  
  comb : process (addr)
  begin
    case conv_integer(addr) is
    when 16#0000# => romdata <= X"88100000";
    when 16#0001# => romdata <= X"0910002B";
    when 16#0002# => romdata <= X"81C12114";
    when 16#0003# => romdata <= X"01000000";
    when 16#0004# => romdata <= X"A1480000";
    when 16#0005# => romdata <= X"A7500000";
    when 16#0006# => romdata <= X"10802B39";
    when 16#0007# => romdata <= X"AC102001";
    when 16#0008# => romdata <= X"91D02000";
    when 16#0009# => romdata <= X"01000000";
    when 16#000A# => romdata <= X"01000000";
    when 16#000B# => romdata <= X"01000000";
    when 16#000C# => romdata <= X"91D02000";
    when 16#000D# => romdata <= X"01000000";
    when 16#000E# => romdata <= X"01000000";
    when 16#000F# => romdata <= X"01000000";
    when 16#0010# => romdata <= X"A1480000";
    when 16#0011# => romdata <= X"29100029";
    when 16#0012# => romdata <= X"81C52150";
    when 16#0013# => romdata <= X"01000000";
    when 16#0014# => romdata <= X"A1480000";
    when 16#0015# => romdata <= X"29100028";
    when 16#0016# => romdata <= X"81C52254";
    when 16#0017# => romdata <= X"01000000";
    when 16#0018# => romdata <= X"A1480000";
    when 16#0019# => romdata <= X"29100028";
    when 16#001A# => romdata <= X"81C522C0";
    when 16#001B# => romdata <= X"01000000";
    when 16#001C# => romdata <= X"91D02000";
    when 16#001D# => romdata <= X"01000000";
    when 16#001E# => romdata <= X"01000000";
    when 16#001F# => romdata <= X"01000000";
    when 16#0020# => romdata <= X"91D02000";
    when 16#0021# => romdata <= X"01000000";
    when 16#0022# => romdata <= X"01000000";
    when 16#0023# => romdata <= X"01000000";
    when 16#0024# => romdata <= X"A1480000";
    when 16#0025# => romdata <= X"A7500000";
    when 16#0026# => romdata <= X"10802B19";
    when 16#0027# => romdata <= X"AC102009";
    when 16#0028# => romdata <= X"91D02000";
    when 16#0029# => romdata <= X"01000000";
    when 16#002A# => romdata <= X"01000000";
    when 16#002B# => romdata <= X"01000000";
    when 16#002C# => romdata <= X"91D02000";
    when 16#002D# => romdata <= X"01000000";
    when 16#002E# => romdata <= X"01000000";
    when 16#002F# => romdata <= X"01000000";
    when 16#0030# => romdata <= X"91D02000";
    when 16#0031# => romdata <= X"01000000";
    when 16#0032# => romdata <= X"01000000";
    when 16#0033# => romdata <= X"01000000";
    when 16#0034# => romdata <= X"91D02000";
    when 16#0035# => romdata <= X"01000000";
    when 16#0036# => romdata <= X"01000000";
    when 16#0037# => romdata <= X"01000000";
    when 16#0038# => romdata <= X"91D02000";
    when 16#0039# => romdata <= X"01000000";
    when 16#003A# => romdata <= X"01000000";
    when 16#003B# => romdata <= X"01000000";
    when 16#003C# => romdata <= X"91D02000";
    when 16#003D# => romdata <= X"01000000";
    when 16#003E# => romdata <= X"01000000";
    when 16#003F# => romdata <= X"01000000";
    when 16#0040# => romdata <= X"91D02000";
    when 16#0041# => romdata <= X"01000000";
    when 16#0042# => romdata <= X"01000000";
    when 16#0043# => romdata <= X"01000000";
    when 16#0044# => romdata <= X"AE102001";
    when 16#0045# => romdata <= X"A1480000";
    when 16#0046# => romdata <= X"1080295D";
    when 16#0047# => romdata <= X"A7500000";
    when 16#0048# => romdata <= X"AE102002";
    when 16#0049# => romdata <= X"A1480000";
    when 16#004A# => romdata <= X"10802959";
    when 16#004B# => romdata <= X"A7500000";
    when 16#004C# => romdata <= X"AE102003";
    when 16#004D# => romdata <= X"A1480000";
    when 16#004E# => romdata <= X"10802955";
    when 16#004F# => romdata <= X"A7500000";
    when 16#0050# => romdata <= X"AE102004";
    when 16#0051# => romdata <= X"A1480000";
    when 16#0052# => romdata <= X"10802951";
    when 16#0053# => romdata <= X"A7500000";
    when 16#0054# => romdata <= X"AE102005";
    when 16#0055# => romdata <= X"A1480000";
    when 16#0056# => romdata <= X"1080294D";
    when 16#0057# => romdata <= X"A7500000";
    when 16#0058# => romdata <= X"AE102006";
    when 16#0059# => romdata <= X"A1480000";
    when 16#005A# => romdata <= X"10802949";
    when 16#005B# => romdata <= X"A7500000";
    when 16#005C# => romdata <= X"AE102007";
    when 16#005D# => romdata <= X"A1480000";
    when 16#005E# => romdata <= X"10802945";
    when 16#005F# => romdata <= X"A7500000";
    when 16#0060# => romdata <= X"AE102008";
    when 16#0061# => romdata <= X"A1480000";
    when 16#0062# => romdata <= X"10802941";
    when 16#0063# => romdata <= X"A7500000";
    when 16#0064# => romdata <= X"AE102009";
    when 16#0065# => romdata <= X"A1480000";
    when 16#0066# => romdata <= X"1080293D";
    when 16#0067# => romdata <= X"A7500000";
    when 16#0068# => romdata <= X"AE10200A";
    when 16#0069# => romdata <= X"A1480000";
    when 16#006A# => romdata <= X"10802939";
    when 16#006B# => romdata <= X"A7500000";
    when 16#006C# => romdata <= X"AE10200B";
    when 16#006D# => romdata <= X"A1480000";
    when 16#006E# => romdata <= X"10802935";
    when 16#006F# => romdata <= X"A7500000";
    when 16#0070# => romdata <= X"AE10200C";
    when 16#0071# => romdata <= X"A1480000";
    when 16#0072# => romdata <= X"10802931";
    when 16#0073# => romdata <= X"A7500000";
    when 16#0074# => romdata <= X"AE10200D";
    when 16#0075# => romdata <= X"A1480000";
    when 16#0076# => romdata <= X"1080292D";
    when 16#0077# => romdata <= X"A7500000";
    when 16#0078# => romdata <= X"AE10200E";
    when 16#0079# => romdata <= X"A1480000";
    when 16#007A# => romdata <= X"10802929";
    when 16#007B# => romdata <= X"A7500000";
    when 16#007C# => romdata <= X"AE10200F";
    when 16#007D# => romdata <= X"A1480000";
    when 16#007E# => romdata <= X"10802925";
    when 16#007F# => romdata <= X"A7500000";
    when 16#0080# => romdata <= X"91D02000";
    when 16#0081# => romdata <= X"01000000";
    when 16#0082# => romdata <= X"01000000";
    when 16#0083# => romdata <= X"01000000";
    when 16#0084# => romdata <= X"91D02000";
    when 16#0085# => romdata <= X"01000000";
    when 16#0086# => romdata <= X"01000000";
    when 16#0087# => romdata <= X"01000000";
    when 16#0088# => romdata <= X"91D02000";
    when 16#0089# => romdata <= X"01000000";
    when 16#008A# => romdata <= X"01000000";
    when 16#008B# => romdata <= X"01000000";
    when 16#008C# => romdata <= X"91D02000";
    when 16#008D# => romdata <= X"01000000";
    when 16#008E# => romdata <= X"01000000";
    when 16#008F# => romdata <= X"01000000";
    when 16#0090# => romdata <= X"91D02000";
    when 16#0091# => romdata <= X"01000000";
    when 16#0092# => romdata <= X"01000000";
    when 16#0093# => romdata <= X"01000000";
    when 16#0094# => romdata <= X"91D02000";
    when 16#0095# => romdata <= X"01000000";
    when 16#0096# => romdata <= X"01000000";
    when 16#0097# => romdata <= X"01000000";
    when 16#0098# => romdata <= X"91D02000";
    when 16#0099# => romdata <= X"01000000";
    when 16#009A# => romdata <= X"01000000";
    when 16#009B# => romdata <= X"01000000";
    when 16#009C# => romdata <= X"91D02000";
    when 16#009D# => romdata <= X"01000000";
    when 16#009E# => romdata <= X"01000000";
    when 16#009F# => romdata <= X"01000000";
    when 16#00A0# => romdata <= X"91D02000";
    when 16#00A1# => romdata <= X"01000000";
    when 16#00A2# => romdata <= X"01000000";
    when 16#00A3# => romdata <= X"01000000";
    when 16#00A4# => romdata <= X"91D02000";
    when 16#00A5# => romdata <= X"01000000";
    when 16#00A6# => romdata <= X"01000000";
    when 16#00A7# => romdata <= X"01000000";
    when 16#00A8# => romdata <= X"91D02000";
    when 16#00A9# => romdata <= X"01000000";
    when 16#00AA# => romdata <= X"01000000";
    when 16#00AB# => romdata <= X"01000000";
    when 16#00AC# => romdata <= X"91D02000";
    when 16#00AD# => romdata <= X"01000000";
    when 16#00AE# => romdata <= X"01000000";
    when 16#00AF# => romdata <= X"01000000";
    when 16#00B0# => romdata <= X"91D02000";
    when 16#00B1# => romdata <= X"01000000";
    when 16#00B2# => romdata <= X"01000000";
    when 16#00B3# => romdata <= X"01000000";
    when 16#00B4# => romdata <= X"91D02000";
    when 16#00B5# => romdata <= X"01000000";
    when 16#00B6# => romdata <= X"01000000";
    when 16#00B7# => romdata <= X"01000000";
    when 16#00B8# => romdata <= X"91D02000";
    when 16#00B9# => romdata <= X"01000000";
    when 16#00BA# => romdata <= X"01000000";
    when 16#00BB# => romdata <= X"01000000";
    when 16#00BC# => romdata <= X"91D02000";
    when 16#00BD# => romdata <= X"01000000";
    when 16#00BE# => romdata <= X"01000000";
    when 16#00BF# => romdata <= X"01000000";
    when 16#00C0# => romdata <= X"91D02000";
    when 16#00C1# => romdata <= X"01000000";
    when 16#00C2# => romdata <= X"01000000";
    when 16#00C3# => romdata <= X"01000000";
    when 16#00C4# => romdata <= X"91D02000";
    when 16#00C5# => romdata <= X"01000000";
    when 16#00C6# => romdata <= X"01000000";
    when 16#00C7# => romdata <= X"01000000";
    when 16#00C8# => romdata <= X"91D02000";
    when 16#00C9# => romdata <= X"01000000";
    when 16#00CA# => romdata <= X"01000000";
    when 16#00CB# => romdata <= X"01000000";
    when 16#00CC# => romdata <= X"91D02000";
    when 16#00CD# => romdata <= X"01000000";
    when 16#00CE# => romdata <= X"01000000";
    when 16#00CF# => romdata <= X"01000000";
    when 16#00D0# => romdata <= X"91D02000";
    when 16#00D1# => romdata <= X"01000000";
    when 16#00D2# => romdata <= X"01000000";
    when 16#00D3# => romdata <= X"01000000";
    when 16#00D4# => romdata <= X"91D02000";
    when 16#00D5# => romdata <= X"01000000";
    when 16#00D6# => romdata <= X"01000000";
    when 16#00D7# => romdata <= X"01000000";
    when 16#00D8# => romdata <= X"91D02000";
    when 16#00D9# => romdata <= X"01000000";
    when 16#00DA# => romdata <= X"01000000";
    when 16#00DB# => romdata <= X"01000000";
    when 16#00DC# => romdata <= X"91D02000";
    when 16#00DD# => romdata <= X"01000000";
    when 16#00DE# => romdata <= X"01000000";
    when 16#00DF# => romdata <= X"01000000";
    when 16#00E0# => romdata <= X"91D02000";
    when 16#00E1# => romdata <= X"01000000";
    when 16#00E2# => romdata <= X"01000000";
    when 16#00E3# => romdata <= X"01000000";
    when 16#00E4# => romdata <= X"91D02000";
    when 16#00E5# => romdata <= X"01000000";
    when 16#00E6# => romdata <= X"01000000";
    when 16#00E7# => romdata <= X"01000000";
    when 16#00E8# => romdata <= X"91D02000";
    when 16#00E9# => romdata <= X"01000000";
    when 16#00EA# => romdata <= X"01000000";
    when 16#00EB# => romdata <= X"01000000";
    when 16#00EC# => romdata <= X"91D02000";
    when 16#00ED# => romdata <= X"01000000";
    when 16#00EE# => romdata <= X"01000000";
    when 16#00EF# => romdata <= X"01000000";
    when 16#00F0# => romdata <= X"91D02000";
    when 16#00F1# => romdata <= X"01000000";
    when 16#00F2# => romdata <= X"01000000";
    when 16#00F3# => romdata <= X"01000000";
    when 16#00F4# => romdata <= X"91D02000";
    when 16#00F5# => romdata <= X"01000000";
    when 16#00F6# => romdata <= X"01000000";
    when 16#00F7# => romdata <= X"01000000";
    when 16#00F8# => romdata <= X"91D02000";
    when 16#00F9# => romdata <= X"01000000";
    when 16#00FA# => romdata <= X"01000000";
    when 16#00FB# => romdata <= X"01000000";
    when 16#00FC# => romdata <= X"91D02000";
    when 16#00FD# => romdata <= X"01000000";
    when 16#00FE# => romdata <= X"01000000";
    when 16#00FF# => romdata <= X"01000000";
    when 16#0100# => romdata <= X"91D02000";
    when 16#0101# => romdata <= X"01000000";
    when 16#0102# => romdata <= X"01000000";
    when 16#0103# => romdata <= X"01000000";
    when 16#0104# => romdata <= X"91D02000";
    when 16#0105# => romdata <= X"01000000";
    when 16#0106# => romdata <= X"01000000";
    when 16#0107# => romdata <= X"01000000";
    when 16#0108# => romdata <= X"91D02000";
    when 16#0109# => romdata <= X"01000000";
    when 16#010A# => romdata <= X"01000000";
    when 16#010B# => romdata <= X"01000000";
    when 16#010C# => romdata <= X"91D02000";
    when 16#010D# => romdata <= X"01000000";
    when 16#010E# => romdata <= X"01000000";
    when 16#010F# => romdata <= X"01000000";
    when 16#0110# => romdata <= X"91D02000";
    when 16#0111# => romdata <= X"01000000";
    when 16#0112# => romdata <= X"01000000";
    when 16#0113# => romdata <= X"01000000";
    when 16#0114# => romdata <= X"91D02000";
    when 16#0115# => romdata <= X"01000000";
    when 16#0116# => romdata <= X"01000000";
    when 16#0117# => romdata <= X"01000000";
    when 16#0118# => romdata <= X"91D02000";
    when 16#0119# => romdata <= X"01000000";
    when 16#011A# => romdata <= X"01000000";
    when 16#011B# => romdata <= X"01000000";
    when 16#011C# => romdata <= X"91D02000";
    when 16#011D# => romdata <= X"01000000";
    when 16#011E# => romdata <= X"01000000";
    when 16#011F# => romdata <= X"01000000";
    when 16#0120# => romdata <= X"91D02000";
    when 16#0121# => romdata <= X"01000000";
    when 16#0122# => romdata <= X"01000000";
    when 16#0123# => romdata <= X"01000000";
    when 16#0124# => romdata <= X"91D02000";
    when 16#0125# => romdata <= X"01000000";
    when 16#0126# => romdata <= X"01000000";
    when 16#0127# => romdata <= X"01000000";
    when 16#0128# => romdata <= X"91D02000";
    when 16#0129# => romdata <= X"01000000";
    when 16#012A# => romdata <= X"01000000";
    when 16#012B# => romdata <= X"01000000";
    when 16#012C# => romdata <= X"91D02000";
    when 16#012D# => romdata <= X"01000000";
    when 16#012E# => romdata <= X"01000000";
    when 16#012F# => romdata <= X"01000000";
    when 16#0130# => romdata <= X"91D02000";
    when 16#0131# => romdata <= X"01000000";
    when 16#0132# => romdata <= X"01000000";
    when 16#0133# => romdata <= X"01000000";
    when 16#0134# => romdata <= X"91D02000";
    when 16#0135# => romdata <= X"01000000";
    when 16#0136# => romdata <= X"01000000";
    when 16#0137# => romdata <= X"01000000";
    when 16#0138# => romdata <= X"91D02000";
    when 16#0139# => romdata <= X"01000000";
    when 16#013A# => romdata <= X"01000000";
    when 16#013B# => romdata <= X"01000000";
    when 16#013C# => romdata <= X"91D02000";
    when 16#013D# => romdata <= X"01000000";
    when 16#013E# => romdata <= X"01000000";
    when 16#013F# => romdata <= X"01000000";
    when 16#0140# => romdata <= X"91D02000";
    when 16#0141# => romdata <= X"01000000";
    when 16#0142# => romdata <= X"01000000";
    when 16#0143# => romdata <= X"01000000";
    when 16#0144# => romdata <= X"91D02000";
    when 16#0145# => romdata <= X"01000000";
    when 16#0146# => romdata <= X"01000000";
    when 16#0147# => romdata <= X"01000000";
    when 16#0148# => romdata <= X"91D02000";
    when 16#0149# => romdata <= X"01000000";
    when 16#014A# => romdata <= X"01000000";
    when 16#014B# => romdata <= X"01000000";
    when 16#014C# => romdata <= X"91D02000";
    when 16#014D# => romdata <= X"01000000";
    when 16#014E# => romdata <= X"01000000";
    when 16#014F# => romdata <= X"01000000";
    when 16#0150# => romdata <= X"91D02000";
    when 16#0151# => romdata <= X"01000000";
    when 16#0152# => romdata <= X"01000000";
    when 16#0153# => romdata <= X"01000000";
    when 16#0154# => romdata <= X"91D02000";
    when 16#0155# => romdata <= X"01000000";
    when 16#0156# => romdata <= X"01000000";
    when 16#0157# => romdata <= X"01000000";
    when 16#0158# => romdata <= X"91D02000";
    when 16#0159# => romdata <= X"01000000";
    when 16#015A# => romdata <= X"01000000";
    when 16#015B# => romdata <= X"01000000";
    when 16#015C# => romdata <= X"91D02000";
    when 16#015D# => romdata <= X"01000000";
    when 16#015E# => romdata <= X"01000000";
    when 16#015F# => romdata <= X"01000000";
    when 16#0160# => romdata <= X"91D02000";
    when 16#0161# => romdata <= X"01000000";
    when 16#0162# => romdata <= X"01000000";
    when 16#0163# => romdata <= X"01000000";
    when 16#0164# => romdata <= X"91D02000";
    when 16#0165# => romdata <= X"01000000";
    when 16#0166# => romdata <= X"01000000";
    when 16#0167# => romdata <= X"01000000";
    when 16#0168# => romdata <= X"91D02000";
    when 16#0169# => romdata <= X"01000000";
    when 16#016A# => romdata <= X"01000000";
    when 16#016B# => romdata <= X"01000000";
    when 16#016C# => romdata <= X"91D02000";
    when 16#016D# => romdata <= X"01000000";
    when 16#016E# => romdata <= X"01000000";
    when 16#016F# => romdata <= X"01000000";
    when 16#0170# => romdata <= X"91D02000";
    when 16#0171# => romdata <= X"01000000";
    when 16#0172# => romdata <= X"01000000";
    when 16#0173# => romdata <= X"01000000";
    when 16#0174# => romdata <= X"91D02000";
    when 16#0175# => romdata <= X"01000000";
    when 16#0176# => romdata <= X"01000000";
    when 16#0177# => romdata <= X"01000000";
    when 16#0178# => romdata <= X"91D02000";
    when 16#0179# => romdata <= X"01000000";
    when 16#017A# => romdata <= X"01000000";
    when 16#017B# => romdata <= X"01000000";
    when 16#017C# => romdata <= X"91D02000";
    when 16#017D# => romdata <= X"01000000";
    when 16#017E# => romdata <= X"01000000";
    when 16#017F# => romdata <= X"01000000";
    when 16#0180# => romdata <= X"91D02000";
    when 16#0181# => romdata <= X"01000000";
    when 16#0182# => romdata <= X"01000000";
    when 16#0183# => romdata <= X"01000000";
    when 16#0184# => romdata <= X"91D02000";
    when 16#0185# => romdata <= X"01000000";
    when 16#0186# => romdata <= X"01000000";
    when 16#0187# => romdata <= X"01000000";
    when 16#0188# => romdata <= X"91D02000";
    when 16#0189# => romdata <= X"01000000";
    when 16#018A# => romdata <= X"01000000";
    when 16#018B# => romdata <= X"01000000";
    when 16#018C# => romdata <= X"91D02000";
    when 16#018D# => romdata <= X"01000000";
    when 16#018E# => romdata <= X"01000000";
    when 16#018F# => romdata <= X"01000000";
    when 16#0190# => romdata <= X"91D02000";
    when 16#0191# => romdata <= X"01000000";
    when 16#0192# => romdata <= X"01000000";
    when 16#0193# => romdata <= X"01000000";
    when 16#0194# => romdata <= X"91D02000";
    when 16#0195# => romdata <= X"01000000";
    when 16#0196# => romdata <= X"01000000";
    when 16#0197# => romdata <= X"01000000";
    when 16#0198# => romdata <= X"91D02000";
    when 16#0199# => romdata <= X"01000000";
    when 16#019A# => romdata <= X"01000000";
    when 16#019B# => romdata <= X"01000000";
    when 16#019C# => romdata <= X"91D02000";
    when 16#019D# => romdata <= X"01000000";
    when 16#019E# => romdata <= X"01000000";
    when 16#019F# => romdata <= X"01000000";
    when 16#01A0# => romdata <= X"91D02000";
    when 16#01A1# => romdata <= X"01000000";
    when 16#01A2# => romdata <= X"01000000";
    when 16#01A3# => romdata <= X"01000000";
    when 16#01A4# => romdata <= X"91D02000";
    when 16#01A5# => romdata <= X"01000000";
    when 16#01A6# => romdata <= X"01000000";
    when 16#01A7# => romdata <= X"01000000";
    when 16#01A8# => romdata <= X"91D02000";
    when 16#01A9# => romdata <= X"01000000";
    when 16#01AA# => romdata <= X"01000000";
    when 16#01AB# => romdata <= X"01000000";
    when 16#01AC# => romdata <= X"91D02000";
    when 16#01AD# => romdata <= X"01000000";
    when 16#01AE# => romdata <= X"01000000";
    when 16#01AF# => romdata <= X"01000000";
    when 16#01B0# => romdata <= X"91D02000";
    when 16#01B1# => romdata <= X"01000000";
    when 16#01B2# => romdata <= X"01000000";
    when 16#01B3# => romdata <= X"01000000";
    when 16#01B4# => romdata <= X"91D02000";
    when 16#01B5# => romdata <= X"01000000";
    when 16#01B6# => romdata <= X"01000000";
    when 16#01B7# => romdata <= X"01000000";
    when 16#01B8# => romdata <= X"91D02000";
    when 16#01B9# => romdata <= X"01000000";
    when 16#01BA# => romdata <= X"01000000";
    when 16#01BB# => romdata <= X"01000000";
    when 16#01BC# => romdata <= X"91D02000";
    when 16#01BD# => romdata <= X"01000000";
    when 16#01BE# => romdata <= X"01000000";
    when 16#01BF# => romdata <= X"01000000";
    when 16#01C0# => romdata <= X"91D02000";
    when 16#01C1# => romdata <= X"01000000";
    when 16#01C2# => romdata <= X"01000000";
    when 16#01C3# => romdata <= X"01000000";
    when 16#01C4# => romdata <= X"91D02000";
    when 16#01C5# => romdata <= X"01000000";
    when 16#01C6# => romdata <= X"01000000";
    when 16#01C7# => romdata <= X"01000000";
    when 16#01C8# => romdata <= X"91D02000";
    when 16#01C9# => romdata <= X"01000000";
    when 16#01CA# => romdata <= X"01000000";
    when 16#01CB# => romdata <= X"01000000";
    when 16#01CC# => romdata <= X"91D02000";
    when 16#01CD# => romdata <= X"01000000";
    when 16#01CE# => romdata <= X"01000000";
    when 16#01CF# => romdata <= X"01000000";
    when 16#01D0# => romdata <= X"91D02000";
    when 16#01D1# => romdata <= X"01000000";
    when 16#01D2# => romdata <= X"01000000";
    when 16#01D3# => romdata <= X"01000000";
    when 16#01D4# => romdata <= X"91D02000";
    when 16#01D5# => romdata <= X"01000000";
    when 16#01D6# => romdata <= X"01000000";
    when 16#01D7# => romdata <= X"01000000";
    when 16#01D8# => romdata <= X"91D02000";
    when 16#01D9# => romdata <= X"01000000";
    when 16#01DA# => romdata <= X"01000000";
    when 16#01DB# => romdata <= X"01000000";
    when 16#01DC# => romdata <= X"91D02000";
    when 16#01DD# => romdata <= X"01000000";
    when 16#01DE# => romdata <= X"01000000";
    when 16#01DF# => romdata <= X"01000000";
    when 16#01E0# => romdata <= X"91D02000";
    when 16#01E1# => romdata <= X"01000000";
    when 16#01E2# => romdata <= X"01000000";
    when 16#01E3# => romdata <= X"01000000";
    when 16#01E4# => romdata <= X"91D02000";
    when 16#01E5# => romdata <= X"01000000";
    when 16#01E6# => romdata <= X"01000000";
    when 16#01E7# => romdata <= X"01000000";
    when 16#01E8# => romdata <= X"91D02000";
    when 16#01E9# => romdata <= X"01000000";
    when 16#01EA# => romdata <= X"01000000";
    when 16#01EB# => romdata <= X"01000000";
    when 16#01EC# => romdata <= X"91D02000";
    when 16#01ED# => romdata <= X"01000000";
    when 16#01EE# => romdata <= X"01000000";
    when 16#01EF# => romdata <= X"01000000";
    when 16#01F0# => romdata <= X"91D02000";
    when 16#01F1# => romdata <= X"01000000";
    when 16#01F2# => romdata <= X"01000000";
    when 16#01F3# => romdata <= X"01000000";
    when 16#01F4# => romdata <= X"91D02000";
    when 16#01F5# => romdata <= X"01000000";
    when 16#01F6# => romdata <= X"01000000";
    when 16#01F7# => romdata <= X"01000000";
    when 16#01F8# => romdata <= X"91D02000";
    when 16#01F9# => romdata <= X"01000000";
    when 16#01FA# => romdata <= X"01000000";
    when 16#01FB# => romdata <= X"01000000";
    when 16#01FC# => romdata <= X"91D02000";
    when 16#01FD# => romdata <= X"01000000";
    when 16#01FE# => romdata <= X"01000000";
    when 16#01FF# => romdata <= X"01000000";
    when 16#0200# => romdata <= X"91D02000";
    when 16#0201# => romdata <= X"01000000";
    when 16#0202# => romdata <= X"01000000";
    when 16#0203# => romdata <= X"01000000";
    when 16#0204# => romdata <= X"91D02000";
    when 16#0205# => romdata <= X"01000000";
    when 16#0206# => romdata <= X"01000000";
    when 16#0207# => romdata <= X"01000000";
    when 16#0208# => romdata <= X"A1480000";
    when 16#0209# => romdata <= X"29100029";
    when 16#020A# => romdata <= X"81C52094";
    when 16#020B# => romdata <= X"01000000";
    when 16#020C# => romdata <= X"A1480000";
    when 16#020D# => romdata <= X"108026BC";
    when 16#020E# => romdata <= X"A7500000";
    when 16#020F# => romdata <= X"01000000";
    when 16#0210# => romdata <= X"91D02000";
    when 16#0211# => romdata <= X"01000000";
    when 16#0212# => romdata <= X"01000000";
    when 16#0213# => romdata <= X"01000000";
    when 16#0214# => romdata <= X"A1480000";
    when 16#0215# => romdata <= X"29100029";
    when 16#0216# => romdata <= X"81C52078";
    when 16#0217# => romdata <= X"01000000";
    when 16#0218# => romdata <= X"91D02000";
    when 16#0219# => romdata <= X"01000000";
    when 16#021A# => romdata <= X"01000000";
    when 16#021B# => romdata <= X"01000000";
    when 16#021C# => romdata <= X"91D02000";
    when 16#021D# => romdata <= X"01000000";
    when 16#021E# => romdata <= X"01000000";
    when 16#021F# => romdata <= X"01000000";
    when 16#0220# => romdata <= X"91D02000";
    when 16#0221# => romdata <= X"01000000";
    when 16#0222# => romdata <= X"01000000";
    when 16#0223# => romdata <= X"01000000";
    when 16#0224# => romdata <= X"91D02000";
    when 16#0225# => romdata <= X"01000000";
    when 16#0226# => romdata <= X"01000000";
    when 16#0227# => romdata <= X"01000000";
    when 16#0228# => romdata <= X"91D02000";
    when 16#0229# => romdata <= X"01000000";
    when 16#022A# => romdata <= X"01000000";
    when 16#022B# => romdata <= X"01000000";
    when 16#022C# => romdata <= X"91D02000";
    when 16#022D# => romdata <= X"01000000";
    when 16#022E# => romdata <= X"01000000";
    when 16#022F# => romdata <= X"01000000";
    when 16#0230# => romdata <= X"91D02000";
    when 16#0231# => romdata <= X"01000000";
    when 16#0232# => romdata <= X"01000000";
    when 16#0233# => romdata <= X"01000000";
    when 16#0234# => romdata <= X"91D02000";
    when 16#0235# => romdata <= X"01000000";
    when 16#0236# => romdata <= X"01000000";
    when 16#0237# => romdata <= X"01000000";
    when 16#0238# => romdata <= X"91D02000";
    when 16#0239# => romdata <= X"01000000";
    when 16#023A# => romdata <= X"01000000";
    when 16#023B# => romdata <= X"01000000";
    when 16#023C# => romdata <= X"91D02000";
    when 16#023D# => romdata <= X"01000000";
    when 16#023E# => romdata <= X"01000000";
    when 16#023F# => romdata <= X"01000000";
    when 16#0240# => romdata <= X"91D02000";
    when 16#0241# => romdata <= X"01000000";
    when 16#0242# => romdata <= X"01000000";
    when 16#0243# => romdata <= X"01000000";
    when 16#0244# => romdata <= X"91D02000";
    when 16#0245# => romdata <= X"01000000";
    when 16#0246# => romdata <= X"01000000";
    when 16#0247# => romdata <= X"01000000";
    when 16#0248# => romdata <= X"91D02000";
    when 16#0249# => romdata <= X"01000000";
    when 16#024A# => romdata <= X"01000000";
    when 16#024B# => romdata <= X"01000000";
    when 16#024C# => romdata <= X"91D02000";
    when 16#024D# => romdata <= X"01000000";
    when 16#024E# => romdata <= X"01000000";
    when 16#024F# => romdata <= X"01000000";
    when 16#0250# => romdata <= X"91D02000";
    when 16#0251# => romdata <= X"01000000";
    when 16#0252# => romdata <= X"01000000";
    when 16#0253# => romdata <= X"01000000";
    when 16#0254# => romdata <= X"91D02000";
    when 16#0255# => romdata <= X"01000000";
    when 16#0256# => romdata <= X"01000000";
    when 16#0257# => romdata <= X"01000000";
    when 16#0258# => romdata <= X"91D02000";
    when 16#0259# => romdata <= X"01000000";
    when 16#025A# => romdata <= X"01000000";
    when 16#025B# => romdata <= X"01000000";
    when 16#025C# => romdata <= X"91D02000";
    when 16#025D# => romdata <= X"01000000";
    when 16#025E# => romdata <= X"01000000";
    when 16#025F# => romdata <= X"01000000";
    when 16#0260# => romdata <= X"91D02000";
    when 16#0261# => romdata <= X"01000000";
    when 16#0262# => romdata <= X"01000000";
    when 16#0263# => romdata <= X"01000000";
    when 16#0264# => romdata <= X"91D02000";
    when 16#0265# => romdata <= X"01000000";
    when 16#0266# => romdata <= X"01000000";
    when 16#0267# => romdata <= X"01000000";
    when 16#0268# => romdata <= X"91D02000";
    when 16#0269# => romdata <= X"01000000";
    when 16#026A# => romdata <= X"01000000";
    when 16#026B# => romdata <= X"01000000";
    when 16#026C# => romdata <= X"91D02000";
    when 16#026D# => romdata <= X"01000000";
    when 16#026E# => romdata <= X"01000000";
    when 16#026F# => romdata <= X"01000000";
    when 16#0270# => romdata <= X"91D02000";
    when 16#0271# => romdata <= X"01000000";
    when 16#0272# => romdata <= X"01000000";
    when 16#0273# => romdata <= X"01000000";
    when 16#0274# => romdata <= X"91D02000";
    when 16#0275# => romdata <= X"01000000";
    when 16#0276# => romdata <= X"01000000";
    when 16#0277# => romdata <= X"01000000";
    when 16#0278# => romdata <= X"91D02000";
    when 16#0279# => romdata <= X"01000000";
    when 16#027A# => romdata <= X"01000000";
    when 16#027B# => romdata <= X"01000000";
    when 16#027C# => romdata <= X"91D02000";
    when 16#027D# => romdata <= X"01000000";
    when 16#027E# => romdata <= X"01000000";
    when 16#027F# => romdata <= X"01000000";
    when 16#0280# => romdata <= X"91D02000";
    when 16#0281# => romdata <= X"01000000";
    when 16#0282# => romdata <= X"01000000";
    when 16#0283# => romdata <= X"01000000";
    when 16#0284# => romdata <= X"91D02000";
    when 16#0285# => romdata <= X"01000000";
    when 16#0286# => romdata <= X"01000000";
    when 16#0287# => romdata <= X"01000000";
    when 16#0288# => romdata <= X"91D02000";
    when 16#0289# => romdata <= X"01000000";
    when 16#028A# => romdata <= X"01000000";
    when 16#028B# => romdata <= X"01000000";
    when 16#028C# => romdata <= X"91D02000";
    when 16#028D# => romdata <= X"01000000";
    when 16#028E# => romdata <= X"01000000";
    when 16#028F# => romdata <= X"01000000";
    when 16#0290# => romdata <= X"91D02000";
    when 16#0291# => romdata <= X"01000000";
    when 16#0292# => romdata <= X"01000000";
    when 16#0293# => romdata <= X"01000000";
    when 16#0294# => romdata <= X"91D02000";
    when 16#0295# => romdata <= X"01000000";
    when 16#0296# => romdata <= X"01000000";
    when 16#0297# => romdata <= X"01000000";
    when 16#0298# => romdata <= X"91D02000";
    when 16#0299# => romdata <= X"01000000";
    when 16#029A# => romdata <= X"01000000";
    when 16#029B# => romdata <= X"01000000";
    when 16#029C# => romdata <= X"91D02000";
    when 16#029D# => romdata <= X"01000000";
    when 16#029E# => romdata <= X"01000000";
    when 16#029F# => romdata <= X"01000000";
    when 16#02A0# => romdata <= X"91D02000";
    when 16#02A1# => romdata <= X"01000000";
    when 16#02A2# => romdata <= X"01000000";
    when 16#02A3# => romdata <= X"01000000";
    when 16#02A4# => romdata <= X"91D02000";
    when 16#02A5# => romdata <= X"01000000";
    when 16#02A6# => romdata <= X"01000000";
    when 16#02A7# => romdata <= X"01000000";
    when 16#02A8# => romdata <= X"91D02000";
    when 16#02A9# => romdata <= X"01000000";
    when 16#02AA# => romdata <= X"01000000";
    when 16#02AB# => romdata <= X"01000000";
    when 16#02AC# => romdata <= X"91D02000";
    when 16#02AD# => romdata <= X"01000000";
    when 16#02AE# => romdata <= X"01000000";
    when 16#02AF# => romdata <= X"01000000";
    when 16#02B0# => romdata <= X"91D02000";
    when 16#02B1# => romdata <= X"01000000";
    when 16#02B2# => romdata <= X"01000000";
    when 16#02B3# => romdata <= X"01000000";
    when 16#02B4# => romdata <= X"91D02000";
    when 16#02B5# => romdata <= X"01000000";
    when 16#02B6# => romdata <= X"01000000";
    when 16#02B7# => romdata <= X"01000000";
    when 16#02B8# => romdata <= X"91D02000";
    when 16#02B9# => romdata <= X"01000000";
    when 16#02BA# => romdata <= X"01000000";
    when 16#02BB# => romdata <= X"01000000";
    when 16#02BC# => romdata <= X"91D02000";
    when 16#02BD# => romdata <= X"01000000";
    when 16#02BE# => romdata <= X"01000000";
    when 16#02BF# => romdata <= X"01000000";
    when 16#02C0# => romdata <= X"91D02000";
    when 16#02C1# => romdata <= X"01000000";
    when 16#02C2# => romdata <= X"01000000";
    when 16#02C3# => romdata <= X"01000000";
    when 16#02C4# => romdata <= X"91D02000";
    when 16#02C5# => romdata <= X"01000000";
    when 16#02C6# => romdata <= X"01000000";
    when 16#02C7# => romdata <= X"01000000";
    when 16#02C8# => romdata <= X"91D02000";
    when 16#02C9# => romdata <= X"01000000";
    when 16#02CA# => romdata <= X"01000000";
    when 16#02CB# => romdata <= X"01000000";
    when 16#02CC# => romdata <= X"91D02000";
    when 16#02CD# => romdata <= X"01000000";
    when 16#02CE# => romdata <= X"01000000";
    when 16#02CF# => romdata <= X"01000000";
    when 16#02D0# => romdata <= X"91D02000";
    when 16#02D1# => romdata <= X"01000000";
    when 16#02D2# => romdata <= X"01000000";
    when 16#02D3# => romdata <= X"01000000";
    when 16#02D4# => romdata <= X"91D02000";
    when 16#02D5# => romdata <= X"01000000";
    when 16#02D6# => romdata <= X"01000000";
    when 16#02D7# => romdata <= X"01000000";
    when 16#02D8# => romdata <= X"91D02000";
    when 16#02D9# => romdata <= X"01000000";
    when 16#02DA# => romdata <= X"01000000";
    when 16#02DB# => romdata <= X"01000000";
    when 16#02DC# => romdata <= X"91D02000";
    when 16#02DD# => romdata <= X"01000000";
    when 16#02DE# => romdata <= X"01000000";
    when 16#02DF# => romdata <= X"01000000";
    when 16#02E0# => romdata <= X"91D02000";
    when 16#02E1# => romdata <= X"01000000";
    when 16#02E2# => romdata <= X"01000000";
    when 16#02E3# => romdata <= X"01000000";
    when 16#02E4# => romdata <= X"91D02000";
    when 16#02E5# => romdata <= X"01000000";
    when 16#02E6# => romdata <= X"01000000";
    when 16#02E7# => romdata <= X"01000000";
    when 16#02E8# => romdata <= X"91D02000";
    when 16#02E9# => romdata <= X"01000000";
    when 16#02EA# => romdata <= X"01000000";
    when 16#02EB# => romdata <= X"01000000";
    when 16#02EC# => romdata <= X"91D02000";
    when 16#02ED# => romdata <= X"01000000";
    when 16#02EE# => romdata <= X"01000000";
    when 16#02EF# => romdata <= X"01000000";
    when 16#02F0# => romdata <= X"91D02000";
    when 16#02F1# => romdata <= X"01000000";
    when 16#02F2# => romdata <= X"01000000";
    when 16#02F3# => romdata <= X"01000000";
    when 16#02F4# => romdata <= X"91D02000";
    when 16#02F5# => romdata <= X"01000000";
    when 16#02F6# => romdata <= X"01000000";
    when 16#02F7# => romdata <= X"01000000";
    when 16#02F8# => romdata <= X"91D02000";
    when 16#02F9# => romdata <= X"01000000";
    when 16#02FA# => romdata <= X"01000000";
    when 16#02FB# => romdata <= X"01000000";
    when 16#02FC# => romdata <= X"91D02000";
    when 16#02FD# => romdata <= X"01000000";
    when 16#02FE# => romdata <= X"01000000";
    when 16#02FF# => romdata <= X"01000000";
    when 16#0300# => romdata <= X"91D02000";
    when 16#0301# => romdata <= X"01000000";
    when 16#0302# => romdata <= X"01000000";
    when 16#0303# => romdata <= X"01000000";
    when 16#0304# => romdata <= X"91D02000";
    when 16#0305# => romdata <= X"01000000";
    when 16#0306# => romdata <= X"01000000";
    when 16#0307# => romdata <= X"01000000";
    when 16#0308# => romdata <= X"91D02000";
    when 16#0309# => romdata <= X"01000000";
    when 16#030A# => romdata <= X"01000000";
    when 16#030B# => romdata <= X"01000000";
    when 16#030C# => romdata <= X"91D02000";
    when 16#030D# => romdata <= X"01000000";
    when 16#030E# => romdata <= X"01000000";
    when 16#030F# => romdata <= X"01000000";
    when 16#0310# => romdata <= X"91D02000";
    when 16#0311# => romdata <= X"01000000";
    when 16#0312# => romdata <= X"01000000";
    when 16#0313# => romdata <= X"01000000";
    when 16#0314# => romdata <= X"91D02000";
    when 16#0315# => romdata <= X"01000000";
    when 16#0316# => romdata <= X"01000000";
    when 16#0317# => romdata <= X"01000000";
    when 16#0318# => romdata <= X"91D02000";
    when 16#0319# => romdata <= X"01000000";
    when 16#031A# => romdata <= X"01000000";
    when 16#031B# => romdata <= X"01000000";
    when 16#031C# => romdata <= X"91D02000";
    when 16#031D# => romdata <= X"01000000";
    when 16#031E# => romdata <= X"01000000";
    when 16#031F# => romdata <= X"01000000";
    when 16#0320# => romdata <= X"91D02000";
    when 16#0321# => romdata <= X"01000000";
    when 16#0322# => romdata <= X"01000000";
    when 16#0323# => romdata <= X"01000000";
    when 16#0324# => romdata <= X"91D02000";
    when 16#0325# => romdata <= X"01000000";
    when 16#0326# => romdata <= X"01000000";
    when 16#0327# => romdata <= X"01000000";
    when 16#0328# => romdata <= X"91D02000";
    when 16#0329# => romdata <= X"01000000";
    when 16#032A# => romdata <= X"01000000";
    when 16#032B# => romdata <= X"01000000";
    when 16#032C# => romdata <= X"91D02000";
    when 16#032D# => romdata <= X"01000000";
    when 16#032E# => romdata <= X"01000000";
    when 16#032F# => romdata <= X"01000000";
    when 16#0330# => romdata <= X"91D02000";
    when 16#0331# => romdata <= X"01000000";
    when 16#0332# => romdata <= X"01000000";
    when 16#0333# => romdata <= X"01000000";
    when 16#0334# => romdata <= X"91D02000";
    when 16#0335# => romdata <= X"01000000";
    when 16#0336# => romdata <= X"01000000";
    when 16#0337# => romdata <= X"01000000";
    when 16#0338# => romdata <= X"91D02000";
    when 16#0339# => romdata <= X"01000000";
    when 16#033A# => romdata <= X"01000000";
    when 16#033B# => romdata <= X"01000000";
    when 16#033C# => romdata <= X"91D02000";
    when 16#033D# => romdata <= X"01000000";
    when 16#033E# => romdata <= X"01000000";
    when 16#033F# => romdata <= X"01000000";
    when 16#0340# => romdata <= X"91D02000";
    when 16#0341# => romdata <= X"01000000";
    when 16#0342# => romdata <= X"01000000";
    when 16#0343# => romdata <= X"01000000";
    when 16#0344# => romdata <= X"91D02000";
    when 16#0345# => romdata <= X"01000000";
    when 16#0346# => romdata <= X"01000000";
    when 16#0347# => romdata <= X"01000000";
    when 16#0348# => romdata <= X"91D02000";
    when 16#0349# => romdata <= X"01000000";
    when 16#034A# => romdata <= X"01000000";
    when 16#034B# => romdata <= X"01000000";
    when 16#034C# => romdata <= X"91D02000";
    when 16#034D# => romdata <= X"01000000";
    when 16#034E# => romdata <= X"01000000";
    when 16#034F# => romdata <= X"01000000";
    when 16#0350# => romdata <= X"91D02000";
    when 16#0351# => romdata <= X"01000000";
    when 16#0352# => romdata <= X"01000000";
    when 16#0353# => romdata <= X"01000000";
    when 16#0354# => romdata <= X"91D02000";
    when 16#0355# => romdata <= X"01000000";
    when 16#0356# => romdata <= X"01000000";
    when 16#0357# => romdata <= X"01000000";
    when 16#0358# => romdata <= X"91D02000";
    when 16#0359# => romdata <= X"01000000";
    when 16#035A# => romdata <= X"01000000";
    when 16#035B# => romdata <= X"01000000";
    when 16#035C# => romdata <= X"91D02000";
    when 16#035D# => romdata <= X"01000000";
    when 16#035E# => romdata <= X"01000000";
    when 16#035F# => romdata <= X"01000000";
    when 16#0360# => romdata <= X"91D02000";
    when 16#0361# => romdata <= X"01000000";
    when 16#0362# => romdata <= X"01000000";
    when 16#0363# => romdata <= X"01000000";
    when 16#0364# => romdata <= X"91D02000";
    when 16#0365# => romdata <= X"01000000";
    when 16#0366# => romdata <= X"01000000";
    when 16#0367# => romdata <= X"01000000";
    when 16#0368# => romdata <= X"91D02000";
    when 16#0369# => romdata <= X"01000000";
    when 16#036A# => romdata <= X"01000000";
    when 16#036B# => romdata <= X"01000000";
    when 16#036C# => romdata <= X"91D02000";
    when 16#036D# => romdata <= X"01000000";
    when 16#036E# => romdata <= X"01000000";
    when 16#036F# => romdata <= X"01000000";
    when 16#0370# => romdata <= X"91D02000";
    when 16#0371# => romdata <= X"01000000";
    when 16#0372# => romdata <= X"01000000";
    when 16#0373# => romdata <= X"01000000";
    when 16#0374# => romdata <= X"91D02000";
    when 16#0375# => romdata <= X"01000000";
    when 16#0376# => romdata <= X"01000000";
    when 16#0377# => romdata <= X"01000000";
    when 16#0378# => romdata <= X"91D02000";
    when 16#0379# => romdata <= X"01000000";
    when 16#037A# => romdata <= X"01000000";
    when 16#037B# => romdata <= X"01000000";
    when 16#037C# => romdata <= X"91D02000";
    when 16#037D# => romdata <= X"01000000";
    when 16#037E# => romdata <= X"01000000";
    when 16#037F# => romdata <= X"01000000";
    when 16#0380# => romdata <= X"91D02000";
    when 16#0381# => romdata <= X"01000000";
    when 16#0382# => romdata <= X"01000000";
    when 16#0383# => romdata <= X"01000000";
    when 16#0384# => romdata <= X"91D02000";
    when 16#0385# => romdata <= X"01000000";
    when 16#0386# => romdata <= X"01000000";
    when 16#0387# => romdata <= X"01000000";
    when 16#0388# => romdata <= X"91D02000";
    when 16#0389# => romdata <= X"01000000";
    when 16#038A# => romdata <= X"01000000";
    when 16#038B# => romdata <= X"01000000";
    when 16#038C# => romdata <= X"91D02000";
    when 16#038D# => romdata <= X"01000000";
    when 16#038E# => romdata <= X"01000000";
    when 16#038F# => romdata <= X"01000000";
    when 16#0390# => romdata <= X"91D02000";
    when 16#0391# => romdata <= X"01000000";
    when 16#0392# => romdata <= X"01000000";
    when 16#0393# => romdata <= X"01000000";
    when 16#0394# => romdata <= X"91D02000";
    when 16#0395# => romdata <= X"01000000";
    when 16#0396# => romdata <= X"01000000";
    when 16#0397# => romdata <= X"01000000";
    when 16#0398# => romdata <= X"91D02000";
    when 16#0399# => romdata <= X"01000000";
    when 16#039A# => romdata <= X"01000000";
    when 16#039B# => romdata <= X"01000000";
    when 16#039C# => romdata <= X"91D02000";
    when 16#039D# => romdata <= X"01000000";
    when 16#039E# => romdata <= X"01000000";
    when 16#039F# => romdata <= X"01000000";
    when 16#03A0# => romdata <= X"91D02000";
    when 16#03A1# => romdata <= X"01000000";
    when 16#03A2# => romdata <= X"01000000";
    when 16#03A3# => romdata <= X"01000000";
    when 16#03A4# => romdata <= X"91D02000";
    when 16#03A5# => romdata <= X"01000000";
    when 16#03A6# => romdata <= X"01000000";
    when 16#03A7# => romdata <= X"01000000";
    when 16#03A8# => romdata <= X"91D02000";
    when 16#03A9# => romdata <= X"01000000";
    when 16#03AA# => romdata <= X"01000000";
    when 16#03AB# => romdata <= X"01000000";
    when 16#03AC# => romdata <= X"91D02000";
    when 16#03AD# => romdata <= X"01000000";
    when 16#03AE# => romdata <= X"01000000";
    when 16#03AF# => romdata <= X"01000000";
    when 16#03B0# => romdata <= X"91D02000";
    when 16#03B1# => romdata <= X"01000000";
    when 16#03B2# => romdata <= X"01000000";
    when 16#03B3# => romdata <= X"01000000";
    when 16#03B4# => romdata <= X"91D02000";
    when 16#03B5# => romdata <= X"01000000";
    when 16#03B6# => romdata <= X"01000000";
    when 16#03B7# => romdata <= X"01000000";
    when 16#03B8# => romdata <= X"91D02000";
    when 16#03B9# => romdata <= X"01000000";
    when 16#03BA# => romdata <= X"01000000";
    when 16#03BB# => romdata <= X"01000000";
    when 16#03BC# => romdata <= X"91D02000";
    when 16#03BD# => romdata <= X"01000000";
    when 16#03BE# => romdata <= X"01000000";
    when 16#03BF# => romdata <= X"01000000";
    when 16#03C0# => romdata <= X"91D02000";
    when 16#03C1# => romdata <= X"01000000";
    when 16#03C2# => romdata <= X"01000000";
    when 16#03C3# => romdata <= X"01000000";
    when 16#03C4# => romdata <= X"91D02000";
    when 16#03C5# => romdata <= X"01000000";
    when 16#03C6# => romdata <= X"01000000";
    when 16#03C7# => romdata <= X"01000000";
    when 16#03C8# => romdata <= X"91D02000";
    when 16#03C9# => romdata <= X"01000000";
    when 16#03CA# => romdata <= X"01000000";
    when 16#03CB# => romdata <= X"01000000";
    when 16#03CC# => romdata <= X"91D02000";
    when 16#03CD# => romdata <= X"01000000";
    when 16#03CE# => romdata <= X"01000000";
    when 16#03CF# => romdata <= X"01000000";
    when 16#03D0# => romdata <= X"91D02000";
    when 16#03D1# => romdata <= X"01000000";
    when 16#03D2# => romdata <= X"01000000";
    when 16#03D3# => romdata <= X"01000000";
    when 16#03D4# => romdata <= X"91D02000";
    when 16#03D5# => romdata <= X"01000000";
    when 16#03D6# => romdata <= X"01000000";
    when 16#03D7# => romdata <= X"01000000";
    when 16#03D8# => romdata <= X"91D02000";
    when 16#03D9# => romdata <= X"01000000";
    when 16#03DA# => romdata <= X"01000000";
    when 16#03DB# => romdata <= X"01000000";
    when 16#03DC# => romdata <= X"91D02000";
    when 16#03DD# => romdata <= X"01000000";
    when 16#03DE# => romdata <= X"01000000";
    when 16#03DF# => romdata <= X"01000000";
    when 16#03E0# => romdata <= X"91D02000";
    when 16#03E1# => romdata <= X"01000000";
    when 16#03E2# => romdata <= X"01000000";
    when 16#03E3# => romdata <= X"01000000";
    when 16#03E4# => romdata <= X"91D02000";
    when 16#03E5# => romdata <= X"01000000";
    when 16#03E6# => romdata <= X"01000000";
    when 16#03E7# => romdata <= X"01000000";
    when 16#03E8# => romdata <= X"91D02000";
    when 16#03E9# => romdata <= X"01000000";
    when 16#03EA# => romdata <= X"01000000";
    when 16#03EB# => romdata <= X"01000000";
    when 16#03EC# => romdata <= X"91D02000";
    when 16#03ED# => romdata <= X"01000000";
    when 16#03EE# => romdata <= X"01000000";
    when 16#03EF# => romdata <= X"01000000";
    when 16#03F0# => romdata <= X"91D02000";
    when 16#03F1# => romdata <= X"01000000";
    when 16#03F2# => romdata <= X"01000000";
    when 16#03F3# => romdata <= X"01000000";
    when 16#03F4# => romdata <= X"91D02000";
    when 16#03F5# => romdata <= X"01000000";
    when 16#03F6# => romdata <= X"01000000";
    when 16#03F7# => romdata <= X"01000000";
    when 16#03F8# => romdata <= X"91D02000";
    when 16#03F9# => romdata <= X"01000000";
    when 16#03FA# => romdata <= X"01000000";
    when 16#03FB# => romdata <= X"01000000";
    when 16#03FC# => romdata <= X"91D02000";
    when 16#03FD# => romdata <= X"01000000";
    when 16#03FE# => romdata <= X"01000000";
    when 16#03FF# => romdata <= X"01000000";
    when 16#0400# => romdata <= X"9DE3BFC0";
    when 16#0401# => romdata <= X"05100035";
    when 16#0402# => romdata <= X"8410A230";
    when 16#0403# => romdata <= X"07100038";
    when 16#0404# => romdata <= X"8610E278";
    when 16#0405# => romdata <= X"82100000";
    when 16#0406# => romdata <= X"8620C002";
    when 16#0407# => romdata <= X"86A0E008";
    when 16#0408# => romdata <= X"36BFFFFF";
    when 16#0409# => romdata <= X"C0388003";
    when 16#040A# => romdata <= X"11100038";
    when 16#040B# => romdata <= X"90122278";
    when 16#040C# => romdata <= X"C0220000";
    when 16#040D# => romdata <= X"40002590";
    when 16#040E# => romdata <= X"01000000";
    when 16#040F# => romdata <= X"40002590";
    when 16#0410# => romdata <= X"01000000";
    when 16#0411# => romdata <= X"40002742";
    when 16#0412# => romdata <= X"01000000";
    when 16#0413# => romdata <= X"11100032";
    when 16#0414# => romdata <= X"90122294";
    when 16#0415# => romdata <= X"40000547";
    when 16#0416# => romdata <= X"01000000";
    when 16#0417# => romdata <= X"40002E87";
    when 16#0418# => romdata <= X"01000000";
    when 16#0419# => romdata <= X"40000531";
    when 16#041A# => romdata <= X"01000000";
    when 16#041B# => romdata <= X"4000266D";
    when 16#041C# => romdata <= X"01000000";
    when 16#041D# => romdata <= X"81C7E008";
    when 16#041E# => romdata <= X"81E80000";
    when 16#041F# => romdata <= X"9DE3BFA0";
    when 16#0420# => romdata <= X"21100035";
    when 16#0421# => romdata <= X"C20C2230";
    when 16#0422# => romdata <= X"80A06000";
    when 16#0423# => romdata <= X"12800022";
    when 16#0424# => romdata <= X"23100035";
    when 16#0425# => romdata <= X"C2046234";
    when 16#0426# => romdata <= X"27100030";
    when 16#0427# => romdata <= X"25100030";
    when 16#0428# => romdata <= X"A614E0EC";
    when 16#0429# => romdata <= X"A414A0F0";
    when 16#042A# => romdata <= X"A4248013";
    when 16#042B# => romdata <= X"A53CA002";
    when 16#042C# => romdata <= X"A404BFFF";
    when 16#042D# => romdata <= X"80A04012";
    when 16#042E# => romdata <= X"3A80000E";
    when 16#042F# => romdata <= X"03000000";
    when 16#0430# => romdata <= X"A2146234";
    when 16#0431# => romdata <= X"82006001";
    when 16#0432# => romdata <= X"85286002";
    when 16#0433# => romdata <= X"C2244000";
    when 16#0434# => romdata <= X"C204C002";
    when 16#0435# => romdata <= X"9FC04000";
    when 16#0436# => romdata <= X"01000000";
    when 16#0437# => romdata <= X"C2044000";
    when 16#0438# => romdata <= X"80A04012";
    when 16#0439# => romdata <= X"0ABFFFF9";
    when 16#043A# => romdata <= X"82006001";
    when 16#043B# => romdata <= X"03000000";
    when 16#043C# => romdata <= X"82106000";
    when 16#043D# => romdata <= X"80A06000";
    when 16#043E# => romdata <= X"02800006";
    when 16#043F# => romdata <= X"82102001";
    when 16#0440# => romdata <= X"1110002C";
    when 16#0441# => romdata <= X"6FFFFBBF";
    when 16#0442# => romdata <= X"90122260";
    when 16#0443# => romdata <= X"82102001";
    when 16#0444# => romdata <= X"C22C2230";
    when 16#0445# => romdata <= X"81C7E008";
    when 16#0446# => romdata <= X"81E80000";
    when 16#0447# => romdata <= X"9DE3BFA0";
    when 16#0448# => romdata <= X"81C7E008";
    when 16#0449# => romdata <= X"81E80000";
    when 16#044A# => romdata <= X"9DE3BFA0";
    when 16#044B# => romdata <= X"03000000";
    when 16#044C# => romdata <= X"82106000";
    when 16#044D# => romdata <= X"80A06000";
    when 16#044E# => romdata <= X"22800008";
    when 16#044F# => romdata <= X"11100038";
    when 16#0450# => romdata <= X"1110002C";
    when 16#0451# => romdata <= X"13100035";
    when 16#0452# => romdata <= X"90122260";
    when 16#0453# => romdata <= X"6FFFFBAD";
    when 16#0454# => romdata <= X"92126238";
    when 16#0455# => romdata <= X"11100038";
    when 16#0456# => romdata <= X"C2022278";
    when 16#0457# => romdata <= X"80A06000";
    when 16#0458# => romdata <= X"02800009";
    when 16#0459# => romdata <= X"90122278";
    when 16#045A# => romdata <= X"03000000";
    when 16#045B# => romdata <= X"82106000";
    when 16#045C# => romdata <= X"80A06000";
    when 16#045D# => romdata <= X"02800004";
    when 16#045E# => romdata <= X"01000000";
    when 16#045F# => romdata <= X"9FC04000";
    when 16#0460# => romdata <= X"01000000";
    when 16#0461# => romdata <= X"81C7E008";
    when 16#0462# => romdata <= X"81E80000";
    when 16#0463# => romdata <= X"9DE3BFA0";
    when 16#0464# => romdata <= X"81C7E008";
    when 16#0465# => romdata <= X"81E80000";
    when 16#0466# => romdata <= X"81C3E008";
    when 16#0467# => romdata <= X"01000000";
    when 16#0468# => romdata <= X"03100035";
    when 16#0469# => romdata <= X"81C3E008";
    when 16#046A# => romdata <= X"D0206250";
    when 16#046B# => romdata <= X"03100036";
    when 16#046C# => romdata <= X"81C3E008";
    when 16#046D# => romdata <= X"D0006258";
    when 16#046E# => romdata <= X"9DE3BFA0";
    when 16#046F# => romdata <= X"07100036";
    when 16#0470# => romdata <= X"C200E258";
    when 16#0471# => romdata <= X"80A06000";
    when 16#0472# => romdata <= X"02800018";
    when 16#0473# => romdata <= X"03100035";
    when 16#0474# => romdata <= X"8610E258";
    when 16#0475# => romdata <= X"C4006250";
    when 16#0476# => romdata <= X"03100032";
    when 16#0477# => romdata <= X"DA0062C0";
    when 16#0478# => romdata <= X"C200A004";
    when 16#0479# => romdata <= X"80886200";
    when 16#047A# => romdata <= X"12800015";
    when 16#047B# => romdata <= X"01000000";
    when 16#047C# => romdata <= X"C200C000";
    when 16#047D# => romdata <= X"88200001";
    when 16#047E# => romdata <= X"C84B4004";
    when 16#047F# => romdata <= X"C8208000";
    when 16#0480# => romdata <= X"82007FFF";
    when 16#0481# => romdata <= X"80A06000";
    when 16#0482# => romdata <= X"12BFFFF6";
    when 16#0483# => romdata <= X"C220C000";
    when 16#0484# => romdata <= X"C200A008";
    when 16#0485# => romdata <= X"07000010";
    when 16#0486# => romdata <= X"82284003";
    when 16#0487# => romdata <= X"C220A008";
    when 16#0488# => romdata <= X"81C7E008";
    when 16#0489# => romdata <= X"81E80000";
    when 16#048A# => romdata <= X"07000010";
    when 16#048B# => romdata <= X"C2006250";
    when 16#048C# => romdata <= X"C4006008";
    when 16#048D# => romdata <= X"84288003";
    when 16#048E# => romdata <= X"C4206008";
    when 16#048F# => romdata <= X"81C7E008";
    when 16#0490# => romdata <= X"81E80000";
    when 16#0491# => romdata <= X"9DE3BFA0";
    when 16#0492# => romdata <= X"80A66000";
    when 16#0493# => romdata <= X"04800020";
    when 16#0494# => romdata <= X"1F100036";
    when 16#0495# => romdata <= X"05100032";
    when 16#0496# => romdata <= X"19100036";
    when 16#0497# => romdata <= X"8410A2C0";
    when 16#0498# => romdata <= X"98132258";
    when 16#0499# => romdata <= X"9A13E258";
    when 16#049A# => romdata <= X"82102000";
    when 16#049B# => romdata <= X"90100002";
    when 16#049C# => romdata <= X"92033E00";
    when 16#049D# => romdata <= X"9410000D";
    when 16#049E# => romdata <= X"96102200";
    when 16#049F# => romdata <= X"C80E0001";
    when 16#04A0# => romdata <= X"C6008000";
    when 16#04A1# => romdata <= X"C828C000";
    when 16#04A2# => romdata <= X"C828FE00";
    when 16#04A3# => romdata <= X"C8008000";
    when 16#04A4# => romdata <= X"88012001";
    when 16#04A5# => romdata <= X"C8208000";
    when 16#04A6# => romdata <= X"C6034000";
    when 16#04A7# => romdata <= X"80A1000C";
    when 16#04A8# => romdata <= X"0A800003";
    when 16#04A9# => romdata <= X"8600E001";
    when 16#04AA# => romdata <= X"D2220000";
    when 16#04AB# => romdata <= X"80A0E200";
    when 16#04AC# => romdata <= X"04800003";
    when 16#04AD# => romdata <= X"C6234000";
    when 16#04AE# => romdata <= X"D6228000";
    when 16#04AF# => romdata <= X"82006001";
    when 16#04B0# => romdata <= X"80A04019";
    when 16#04B1# => romdata <= X"32BFFFEF";
    when 16#04B2# => romdata <= X"C80E0001";
    when 16#04B3# => romdata <= X"C203E258";
    when 16#04B4# => romdata <= X"80A06000";
    when 16#04B5# => romdata <= X"02800007";
    when 16#04B6# => romdata <= X"03100035";
    when 16#04B7# => romdata <= X"05000010";
    when 16#04B8# => romdata <= X"C2006250";
    when 16#04B9# => romdata <= X"C6006008";
    when 16#04BA# => romdata <= X"8410C002";
    when 16#04BB# => romdata <= X"C4206008";
    when 16#04BC# => romdata <= X"7FFFFFB2";
    when 16#04BD# => romdata <= X"81E80000";
    when 16#04BE# => romdata <= X"01000000";
    when 16#04BF# => romdata <= X"03100035";
    when 16#04C0# => romdata <= X"C2006250";
    when 16#04C1# => romdata <= X"C2006004";
    when 16#04C2# => romdata <= X"8338601A";
    when 16#04C3# => romdata <= X"8208600F";
    when 16#04C4# => romdata <= X"80A00001";
    when 16#04C5# => romdata <= X"81C3E008";
    when 16#04C6# => romdata <= X"90402000";
    when 16#04C7# => romdata <= X"03100035";
    when 16#04C8# => romdata <= X"C2006250";
    when 16#04C9# => romdata <= X"D0004000";
    when 16#04CA# => romdata <= X"81C3E008";
    when 16#04CB# => romdata <= X"01000000";
    when 16#04CC# => romdata <= X"03100035";
    when 16#04CD# => romdata <= X"C4006250";
    when 16#04CE# => romdata <= X"C200A004";
    when 16#04CF# => romdata <= X"8338601A";
    when 16#04D0# => romdata <= X"8088600F";
    when 16#04D1# => romdata <= X"02BFFFFD";
    when 16#04D2# => romdata <= X"01000000";
    when 16#04D3# => romdata <= X"D0008000";
    when 16#04D4# => romdata <= X"81C3E008";
    when 16#04D5# => romdata <= X"01000000";
    when 16#04D6# => romdata <= X"07100035";
    when 16#04D7# => romdata <= X"88102000";
    when 16#04D8# => romdata <= X"8610E250";
    when 16#04D9# => romdata <= X"C400C000";
    when 16#04DA# => romdata <= X"C200A004";
    when 16#04DB# => romdata <= X"8338601A";
    when 16#04DC# => romdata <= X"8088600F";
    when 16#04DD# => romdata <= X"02BFFFFD";
    when 16#04DE# => romdata <= X"01000000";
    when 16#04DF# => romdata <= X"C2008000";
    when 16#04E0# => romdata <= X"C22A0004";
    when 16#04E1# => romdata <= X"83286018";
    when 16#04E2# => romdata <= X"83386018";
    when 16#04E3# => romdata <= X"80A0600A";
    when 16#04E4# => romdata <= X"12BFFFF5";
    when 16#04E5# => romdata <= X"88012001";
    when 16#04E6# => romdata <= X"88013FFF";
    when 16#04E7# => romdata <= X"C02A0004";
    when 16#04E8# => romdata <= X"88020004";
    when 16#04E9# => romdata <= X"C2493FFF";
    when 16#04EA# => romdata <= X"80A0600D";
    when 16#04EB# => romdata <= X"02800004";
    when 16#04EC# => romdata <= X"01000000";
    when 16#04ED# => romdata <= X"81C3E008";
    when 16#04EE# => romdata <= X"01000000";
    when 16#04EF# => romdata <= X"81C3E008";
    when 16#04F0# => romdata <= X"C0293FFF";
    when 16#04F1# => romdata <= X"9DE3BF98";
    when 16#04F2# => romdata <= X"8207A048";
    when 16#04F3# => romdata <= X"92100018";
    when 16#04F4# => romdata <= X"21100036";
    when 16#04F5# => romdata <= X"F227A048";
    when 16#04F6# => romdata <= X"F427A04C";
    when 16#04F7# => romdata <= X"F627A050";
    when 16#04F8# => romdata <= X"F827A054";
    when 16#04F9# => romdata <= X"FA27A058";
    when 16#04FA# => romdata <= X"94100001";
    when 16#04FB# => romdata <= X"C227BFFC";
    when 16#04FC# => romdata <= X"400004BF";
    when 16#04FD# => romdata <= X"90142260";
    when 16#04FE# => romdata <= X"B0100008";
    when 16#04FF# => romdata <= X"90142260";
    when 16#0500# => romdata <= X"7FFFFF91";
    when 16#0501# => romdata <= X"92100018";
    when 16#0502# => romdata <= X"81C7E008";
    when 16#0503# => romdata <= X"81E80000";
    when 16#0504# => romdata <= X"03100036";
    when 16#0505# => romdata <= X"81C3E008";
    when 16#0506# => romdata <= X"D0006360";
    when 16#0507# => romdata <= X"03100036";
    when 16#0508# => romdata <= X"81C3E008";
    when 16#0509# => romdata <= X"C0206360";
    when 16#050A# => romdata <= X"8213C000";
    when 16#050B# => romdata <= X"7FFFFF63";
    when 16#050C# => romdata <= X"9E104000";
    when 16#050D# => romdata <= X"01000000";
    when 16#050E# => romdata <= X"03100036";
    when 16#050F# => romdata <= X"C4006360";
    when 16#0510# => romdata <= X"92100002";
    when 16#0511# => romdata <= X"8400A001";
    when 16#0512# => romdata <= X"11100030";
    when 16#0513# => romdata <= X"C4206360";
    when 16#0514# => romdata <= X"901220F8";
    when 16#0515# => romdata <= X"8213C000";
    when 16#0516# => romdata <= X"7FFFFFDB";
    when 16#0517# => romdata <= X"9E104000";
    when 16#0518# => romdata <= X"01000000";
    when 16#0519# => romdata <= X"03100036";
    when 16#051A# => romdata <= X"C4006360";
    when 16#051B# => romdata <= X"92100002";
    when 16#051C# => romdata <= X"8400A001";
    when 16#051D# => romdata <= X"11100030";
    when 16#051E# => romdata <= X"C4206360";
    when 16#051F# => romdata <= X"90122118";
    when 16#0520# => romdata <= X"8213C000";
    when 16#0521# => romdata <= X"7FFFFFD0";
    when 16#0522# => romdata <= X"9E104000";
    when 16#0523# => romdata <= X"01000000";
    when 16#0524# => romdata <= X"40001700";
    when 16#0525# => romdata <= X"40001740";
    when 16#0526# => romdata <= X"40001534";
    when 16#0527# => romdata <= X"4000177C";
    when 16#0528# => romdata <= X"400017A8";
    when 16#0529# => romdata <= X"40001708";
    when 16#052A# => romdata <= X"400019B0";
    when 16#052B# => romdata <= X"40001904";
    when 16#052C# => romdata <= X"400018A0";
    when 16#052D# => romdata <= X"40001850";
    when 16#052E# => romdata <= X"4000196C";
    when 16#052F# => romdata <= X"C20A0000";
    when 16#0530# => romdata <= X"80A06024";
    when 16#0531# => romdata <= X"22800004";
    when 16#0532# => romdata <= X"C20A2001";
    when 16#0533# => romdata <= X"81C3E008";
    when 16#0534# => romdata <= X"90102000";
    when 16#0535# => romdata <= X"80A06043";
    when 16#0536# => romdata <= X"12BFFFFD";
    when 16#0537# => romdata <= X"01000000";
    when 16#0538# => romdata <= X"C20A2002";
    when 16#0539# => romdata <= X"80A0604D";
    when 16#053A# => romdata <= X"12BFFFF9";
    when 16#053B# => romdata <= X"01000000";
    when 16#053C# => romdata <= X"C20A2003";
    when 16#053D# => romdata <= X"82186044";
    when 16#053E# => romdata <= X"80A00001";
    when 16#053F# => romdata <= X"81C3E008";
    when 16#0540# => romdata <= X"90603FFF";
    when 16#0541# => romdata <= X"9DE3BF98";
    when 16#0542# => romdata <= X"C027BFFC";
    when 16#0543# => romdata <= X"C20E2006";
    when 16#0544# => romdata <= X"80A06005";
    when 16#0545# => romdata <= X"1880007B";
    when 16#0546# => romdata <= X"C6062008";
    when 16#0547# => romdata <= X"83286002";
    when 16#0548# => romdata <= X"05100005";
    when 16#0549# => romdata <= X"8410A090";
    when 16#054A# => romdata <= X"C2008001";
    when 16#054B# => romdata <= X"81C04000";
    when 16#054C# => romdata <= X"01000000";
    when 16#054D# => romdata <= X"82102001";
    when 16#054E# => romdata <= X"C22E2006";
    when 16#054F# => romdata <= X"D806200C";
    when 16#0550# => romdata <= X"82102000";
    when 16#0551# => romdata <= X"80A32000";
    when 16#0552# => romdata <= X"84102000";
    when 16#0553# => romdata <= X"88102001";
    when 16#0554# => romdata <= X"0280000B";
    when 16#0555# => romdata <= X"9E102001";
    when 16#0556# => romdata <= X"88060001";
    when 16#0557# => romdata <= X"DA004003";
    when 16#0558# => romdata <= X"DA212010";
    when 16#0559# => romdata <= X"8400A001";
    when 16#055A# => romdata <= X"80A0800C";
    when 16#055B# => romdata <= X"0ABFFFFB";
    when 16#055C# => romdata <= X"82006004";
    when 16#055D# => romdata <= X"DE0E2006";
    when 16#055E# => romdata <= X"8810000F";
    when 16#055F# => romdata <= X"82102024";
    when 16#0560# => romdata <= X"C22E2048";
    when 16#0561# => romdata <= X"82102043";
    when 16#0562# => romdata <= X"C22E2049";
    when 16#0563# => romdata <= X"8210204D";
    when 16#0564# => romdata <= X"C22E204A";
    when 16#0565# => romdata <= X"82102044";
    when 16#0566# => romdata <= X"C82E0000";
    when 16#0567# => romdata <= X"C22E204B";
    when 16#0568# => romdata <= X"D82E2001";
    when 16#0569# => romdata <= X"DE2E204C";
    when 16#056A# => romdata <= X"D82E204D";
    when 16#056B# => romdata <= X"84100018";
    when 16#056C# => romdata <= X"82102018";
    when 16#056D# => romdata <= X"8930C001";
    when 16#056E# => romdata <= X"C828A04E";
    when 16#056F# => romdata <= X"C828A002";
    when 16#0570# => romdata <= X"82007FF8";
    when 16#0571# => romdata <= X"80A07FF8";
    when 16#0572# => romdata <= X"12BFFFFB";
    when 16#0573# => romdata <= X"8400A001";
    when 16#0574# => romdata <= X"C40E0000";
    when 16#0575# => romdata <= X"C20E2001";
    when 16#0576# => romdata <= X"C60E2003";
    when 16#0577# => romdata <= X"C80E2002";
    when 16#0578# => romdata <= X"8218C001";
    when 16#0579# => romdata <= X"88190002";
    when 16#057A# => romdata <= X"C40E2004";
    when 16#057B# => romdata <= X"88190002";
    when 16#057C# => romdata <= X"C40E2005";
    when 16#057D# => romdata <= X"C82E0000";
    when 16#057E# => romdata <= X"86184002";
    when 16#057F# => romdata <= X"C82E2052";
    when 16#0580# => romdata <= X"832BE018";
    when 16#0581# => romdata <= X"C62E2001";
    when 16#0582# => romdata <= X"83386018";
    when 16#0583# => romdata <= X"C62E2053";
    when 16#0584# => romdata <= X"80A06001";
    when 16#0585# => romdata <= X"84100004";
    when 16#0586# => romdata <= X"82100003";
    when 16#0587# => romdata <= X"90062048";
    when 16#0588# => romdata <= X"12800031";
    when 16#0589# => romdata <= X"9210200C";
    when 16#058A# => romdata <= X"80A32000";
    when 16#058B# => romdata <= X"02800023";
    when 16#058C# => romdata <= X"90100004";
    when 16#058D# => romdata <= X"92100003";
    when 16#058E# => romdata <= X"9610200A";
    when 16#058F# => romdata <= X"94102000";
    when 16#0590# => romdata <= X"8206000B";
    when 16#0591# => romdata <= X"8602E048";
    when 16#0592# => romdata <= X"DA006006";
    when 16#0593# => romdata <= X"86060003";
    when 16#0594# => romdata <= X"84100018";
    when 16#0595# => romdata <= X"82102018";
    when 16#0596# => romdata <= X"89334001";
    when 16#0597# => romdata <= X"C828C000";
    when 16#0598# => romdata <= X"C828A002";
    when 16#0599# => romdata <= X"82007FF8";
    when 16#059A# => romdata <= X"8400A001";
    when 16#059B# => romdata <= X"80A07FF8";
    when 16#059C# => romdata <= X"12BFFFFA";
    when 16#059D# => romdata <= X"8600E001";
    when 16#059E# => romdata <= X"C20E2002";
    when 16#059F# => romdata <= X"9402A001";
    when 16#05A0# => romdata <= X"C40E2004";
    when 16#05A1# => romdata <= X"C60E2005";
    when 16#05A2# => romdata <= X"84188001";
    when 16#05A3# => romdata <= X"9602E004";
    when 16#05A4# => romdata <= X"84188008";
    when 16#05A5# => romdata <= X"C20E2003";
    when 16#05A6# => romdata <= X"80A2800C";
    when 16#05A7# => romdata <= X"8218C001";
    when 16#05A8# => romdata <= X"90100002";
    when 16#05A9# => romdata <= X"82184009";
    when 16#05AA# => romdata <= X"0ABFFFE6";
    when 16#05AB# => romdata <= X"92100001";
    when 16#05AC# => romdata <= X"C22E2001";
    when 16#05AD# => romdata <= X"C42E0000";
    when 16#05AE# => romdata <= X"992B2002";
    when 16#05AF# => romdata <= X"8606000C";
    when 16#05B0# => romdata <= X"C228E053";
    when 16#05B1# => romdata <= X"C428E052";
    when 16#05B2# => romdata <= X"832BE018";
    when 16#05B3# => romdata <= X"90062048";
    when 16#05B4# => romdata <= X"83386018";
    when 16#05B5# => romdata <= X"80A06001";
    when 16#05B6# => romdata <= X"02800003";
    when 16#05B7# => romdata <= X"9203200C";
    when 16#05B8# => romdata <= X"9210200C";
    when 16#05B9# => romdata <= X"7FFFFED8";
    when 16#05BA# => romdata <= X"01000000";
    when 16#05BB# => romdata <= X"7FFFFEB0";
    when 16#05BC# => romdata <= X"01000000";
    when 16#05BD# => romdata <= X"80A22000";
    when 16#05BE# => romdata <= X"12BFFFFD";
    when 16#05BF# => romdata <= X"01000000";
    when 16#05C0# => romdata <= X"81C7E008";
    when 16#05C1# => romdata <= X"91E82001";
    when 16#05C2# => romdata <= X"11100030";
    when 16#05C3# => romdata <= X"C027BFFC";
    when 16#05C4# => romdata <= X"90122158";
    when 16#05C5# => romdata <= X"7FFFFECC";
    when 16#05C6# => romdata <= X"92102008";
    when 16#05C7# => romdata <= X"7FFFFEA4";
    when 16#05C8# => romdata <= X"01000000";
    when 16#05C9# => romdata <= X"80A22000";
    when 16#05CA# => romdata <= X"12BFFFFD";
    when 16#05CB# => romdata <= X"C207BFFC";
    when 16#05CC# => romdata <= X"9FC04000";
    when 16#05CD# => romdata <= X"B0102001";
    when 16#05CE# => romdata <= X"81C7E008";
    when 16#05CF# => romdata <= X"81E80000";
    when 16#05D0# => romdata <= X"C206200C";
    when 16#05D1# => romdata <= X"80A06000";
    when 16#05D2# => romdata <= X"02BFFFEE";
    when 16#05D3# => romdata <= X"82102000";
    when 16#05D4# => romdata <= X"84102000";
    when 16#05D5# => romdata <= X"88060001";
    when 16#05D6# => romdata <= X"C8012010";
    when 16#05D7# => romdata <= X"C8204003";
    when 16#05D8# => romdata <= X"8400A001";
    when 16#05D9# => romdata <= X"C806200C";
    when 16#05DA# => romdata <= X"80A10002";
    when 16#05DB# => romdata <= X"18BFFFFA";
    when 16#05DC# => romdata <= X"82006004";
    when 16#05DD# => romdata <= X"81C7E008";
    when 16#05DE# => romdata <= X"91E82001";
    when 16#05DF# => romdata <= X"11100030";
    when 16#05E0# => romdata <= X"92102011";
    when 16#05E1# => romdata <= X"7FFFFEB0";
    when 16#05E2# => romdata <= X"90122130";
    when 16#05E3# => romdata <= X"7FFFFE88";
    when 16#05E4# => romdata <= X"01000000";
    when 16#05E5# => romdata <= X"80A22000";
    when 16#05E6# => romdata <= X"12BFFFFD";
    when 16#05E7# => romdata <= X"B0102000";
    when 16#05E8# => romdata <= X"81C7E008";
    when 16#05E9# => romdata <= X"81E80000";
    when 16#05EA# => romdata <= X"82102140";
    when 16#05EB# => romdata <= X"11100030";
    when 16#05EC# => romdata <= X"C227BFFC";
    when 16#05ED# => romdata <= X"90122148";
    when 16#05EE# => romdata <= X"7FFFFEA3";
    when 16#05EF# => romdata <= X"9210200A";
    when 16#05F0# => romdata <= X"7FFFFE7B";
    when 16#05F1# => romdata <= X"01000000";
    when 16#05F2# => romdata <= X"80A22000";
    when 16#05F3# => romdata <= X"12BFFFFD";
    when 16#05F4# => romdata <= X"C207BFFC";
    when 16#05F5# => romdata <= X"9FC04000";
    when 16#05F6# => romdata <= X"B0102001";
    when 16#05F7# => romdata <= X"81C7E008";
    when 16#05F8# => romdata <= X"81E80000";
    when 16#05F9# => romdata <= X"9DE3BFA0";
    when 16#05FA# => romdata <= X"9210200E";
    when 16#05FB# => romdata <= X"11100030";
    when 16#05FC# => romdata <= X"7FFFFE95";
    when 16#05FD# => romdata <= X"90122168";
    when 16#05FE# => romdata <= X"7FFFFECE";
    when 16#05FF# => romdata <= X"21100036";
    when 16#0600# => romdata <= X"2B100037";
    when 16#0601# => romdata <= X"D02C2368";
    when 16#0602# => romdata <= X"AA156068";
    when 16#0603# => romdata <= X"A0142368";
    when 16#0604# => romdata <= X"37100030";
    when 16#0605# => romdata <= X"D02C2080";
    when 16#0606# => romdata <= X"AC042100";
    when 16#0607# => romdata <= X"3B100005";
    when 16#0608# => romdata <= X"B4102000";
    when 16#0609# => romdata <= X"B616E178";
    when 16#060A# => romdata <= X"BA1760A8";
    when 16#060B# => romdata <= X"A0042081";
    when 16#060C# => romdata <= X"B8100015";
    when 16#060D# => romdata <= X"80A6A004";
    when 16#060E# => romdata <= X"38800063";
    when 16#060F# => romdata <= X"80A6A005";
    when 16#0610# => romdata <= X"832EA002";
    when 16#0611# => romdata <= X"C2074001";
    when 16#0612# => romdata <= X"81C04000";
    when 16#0613# => romdata <= X"01000000";
    when 16#0614# => romdata <= X"C20C3FFF";
    when 16#0615# => romdata <= X"840CE0FF";
    when 16#0616# => romdata <= X"860860FF";
    when 16#0617# => romdata <= X"80A0C002";
    when 16#0618# => romdata <= X"02800004";
    when 16#0619# => romdata <= X"B4102004";
    when 16#061A# => romdata <= X"82100013";
    when 16#061B# => romdata <= X"B4102000";
    when 16#061C# => romdata <= X"A4100011";
    when 16#061D# => romdata <= X"A6100001";
    when 16#061E# => romdata <= X"7FFFFEAE";
    when 16#061F# => romdata <= X"01000000";
    when 16#0620# => romdata <= X"D02C0000";
    when 16#0621# => romdata <= X"D02C3F80";
    when 16#0622# => romdata <= X"A0042001";
    when 16#0623# => romdata <= X"80A40016";
    when 16#0624# => romdata <= X"3A800002";
    when 16#0625# => romdata <= X"A0043F80";
    when 16#0626# => romdata <= X"10BFFFE7";
    when 16#0627# => romdata <= X"A2100012";
    when 16#0628# => romdata <= X"C40C3FFF";
    when 16#0629# => romdata <= X"8205E004";
    when 16#062A# => romdata <= X"8808A0FF";
    when 16#062B# => romdata <= X"83286002";
    when 16#062C# => romdata <= X"C6054001";
    when 16#062D# => romdata <= X"8728E008";
    when 16#062E# => romdata <= X"86110003";
    when 16#062F# => romdata <= X"C6254001";
    when 16#0630# => romdata <= X"808D2001";
    when 16#0631# => romdata <= X"02800004";
    when 16#0632# => romdata <= X"82188013";
    when 16#0633# => romdata <= X"A2188011";
    when 16#0634# => romdata <= X"82100013";
    when 16#0635# => romdata <= X"A8052001";
    when 16#0636# => romdata <= X"80A52003";
    when 16#0637# => romdata <= X"08800039";
    when 16#0638# => romdata <= X"A6100001";
    when 16#0639# => romdata <= X"AE05E001";
    when 16#063A# => romdata <= X"C407200C";
    when 16#063B# => romdata <= X"80A5C002";
    when 16#063C# => romdata <= X"2A800044";
    when 16#063D# => romdata <= X"8205E004";
    when 16#063E# => romdata <= X"B4102003";
    when 16#063F# => romdata <= X"10BFFFDD";
    when 16#0640# => romdata <= X"A8102000";
    when 16#0641# => romdata <= X"C4056008";
    when 16#0642# => romdata <= X"C20C3FFF";
    when 16#0643# => romdata <= X"8528A008";
    when 16#0644# => romdata <= X"860860FF";
    when 16#0645# => romdata <= X"8410C002";
    when 16#0646# => romdata <= X"808D2001";
    when 16#0647# => romdata <= X"02800037";
    when 16#0648# => romdata <= X"C4256008";
    when 16#0649# => romdata <= X"A2184011";
    when 16#064A# => romdata <= X"A8052001";
    when 16#064B# => romdata <= X"80A52003";
    when 16#064C# => romdata <= X"08800025";
    when 16#064D# => romdata <= X"80A6A005";
    when 16#064E# => romdata <= X"C0272010";
    when 16#064F# => romdata <= X"C207200C";
    when 16#0650# => romdata <= X"80A06000";
    when 16#0651# => romdata <= X"02800006";
    when 16#0652# => romdata <= X"82100013";
    when 16#0653# => romdata <= X"C24F2006";
    when 16#0654# => romdata <= X"80A06001";
    when 16#0655# => romdata <= X"02800044";
    when 16#0656# => romdata <= X"82100013";
    when 16#0657# => romdata <= X"AE102000";
    when 16#0658# => romdata <= X"B4102003";
    when 16#0659# => romdata <= X"10BFFFC3";
    when 16#065A# => romdata <= X"A8102000";
    when 16#065B# => romdata <= X"E40C3FFF";
    when 16#065C# => romdata <= X"820C60FF";
    when 16#065D# => romdata <= X"840CA0FF";
    when 16#065E# => romdata <= X"80A08001";
    when 16#065F# => romdata <= X"12BFFFBC";
    when 16#0660# => romdata <= X"82100013";
    when 16#0661# => romdata <= X"7FFFFEE0";
    when 16#0662# => romdata <= X"90100015";
    when 16#0663# => romdata <= X"92102005";
    when 16#0664# => romdata <= X"A2100008";
    when 16#0665# => romdata <= X"7FFFFE2C";
    when 16#0666# => romdata <= X"9010001B";
    when 16#0667# => romdata <= X"808C60FF";
    when 16#0668# => romdata <= X"12BFFFB6";
    when 16#0669# => romdata <= X"B4102000";
    when 16#066A# => romdata <= X"81C7E008";
    when 16#066B# => romdata <= X"91E82000";
    when 16#066C# => romdata <= X"C20C3FFA";
    when 16#066D# => romdata <= X"80A06024";
    when 16#066E# => romdata <= X"02800016";
    when 16#066F# => romdata <= X"82043FFA";
    when 16#0670# => romdata <= X"80A6A005";
    when 16#0671# => romdata <= X"A4100011";
    when 16#0672# => romdata <= X"12BFFFAB";
    when 16#0673# => romdata <= X"82100013";
    when 16#0674# => romdata <= X"7FFFFECD";
    when 16#0675# => romdata <= X"90100015";
    when 16#0676# => romdata <= X"92102005";
    when 16#0677# => romdata <= X"A2100008";
    when 16#0678# => romdata <= X"7FFFFE19";
    when 16#0679# => romdata <= X"9010001B";
    when 16#067A# => romdata <= X"808C60FF";
    when 16#067B# => romdata <= X"02BFFFEF";
    when 16#067C# => romdata <= X"B4102000";
    when 16#067D# => romdata <= X"30BFFFA1";
    when 16#067E# => romdata <= X"10BFFFCC";
    when 16#067F# => romdata <= X"A6184013";
    when 16#0680# => romdata <= X"A8102000";
    when 16#0681# => romdata <= X"83286002";
    when 16#0682# => romdata <= X"10BFFFEE";
    when 16#0683# => romdata <= X"C0270001";
    when 16#0684# => romdata <= X"C4086001";
    when 16#0685# => romdata <= X"80A0A043";
    when 16#0686# => romdata <= X"12BFFFEB";
    when 16#0687# => romdata <= X"80A6A005";
    when 16#0688# => romdata <= X"C4086002";
    when 16#0689# => romdata <= X"80A0A04D";
    when 16#068A# => romdata <= X"12BFFFE7";
    when 16#068B# => romdata <= X"80A6A005";
    when 16#068C# => romdata <= X"C2086003";
    when 16#068D# => romdata <= X"80A06044";
    when 16#068E# => romdata <= X"12BFFFE3";
    when 16#068F# => romdata <= X"80A6A005";
    when 16#0690# => romdata <= X"C0256008";
    when 16#0691# => romdata <= X"B4102001";
    when 16#0692# => romdata <= X"C20C3FFE";
    when 16#0693# => romdata <= X"A8102000";
    when 16#0694# => romdata <= X"C22D6006";
    when 16#0695# => romdata <= X"E20C3FFF";
    when 16#0696# => romdata <= X"840C60FF";
    when 16#0697# => romdata <= X"10BFFF85";
    when 16#0698# => romdata <= X"C425600C";
    when 16#0699# => romdata <= X"AE102000";
    when 16#069A# => romdata <= X"B4102002";
    when 16#069B# => romdata <= X"10BFFF81";
    when 16#069C# => romdata <= X"A8102000";
    when 16#069D# => romdata <= X"400022B4";
    when 16#069E# => romdata <= X"4000237C";
    when 16#069F# => romdata <= X"40002370";
    when 16#06A0# => romdata <= X"40002364";
    when 16#06A1# => romdata <= X"40002358";
    when 16#06A2# => romdata <= X"4000234C";
    when 16#06A3# => romdata <= X"4000232C";
    when 16#06A4# => romdata <= X"400022F4";
    when 16#06A5# => romdata <= X"81C3E008";
    when 16#06A6# => romdata <= X"D2222084";
    when 16#06A7# => romdata <= X"80A26000";
    when 16#06A8# => romdata <= X"02800007";
    when 16#06A9# => romdata <= X"80A26001";
    when 16#06AA# => romdata <= X"02800006";
    when 16#06AB# => romdata <= X"82102001";
    when 16#06AC# => romdata <= X"80A260F1";
    when 16#06AD# => romdata <= X"02800003";
    when 16#06AE# => romdata <= X"82102002";
    when 16#06AF# => romdata <= X"82102000";
    when 16#06B0# => romdata <= X"83286003";
    when 16#06B1# => romdata <= X"05100031";
    when 16#06B2# => romdata <= X"8410A3E4";
    when 16#06B3# => romdata <= X"82008001";
    when 16#06B4# => romdata <= X"81C3E008";
    when 16#06B5# => romdata <= X"D0006004";
    when 16#06B6# => romdata <= X"80A26000";
    when 16#06B7# => romdata <= X"0280000C";
    when 16#06B8# => romdata <= X"03100031";
    when 16#06B9# => romdata <= X"84102001";
    when 16#06BA# => romdata <= X"82106374";
    when 16#06BB# => romdata <= X"C6004000";
    when 16#06BC# => romdata <= X"80A0C009";
    when 16#06BD# => romdata <= X"22800008";
    when 16#06BE# => romdata <= X"8528A003";
    when 16#06BF# => romdata <= X"8400A001";
    when 16#06C0# => romdata <= X"80A0A00F";
    when 16#06C1# => romdata <= X"12BFFFFA";
    when 16#06C2# => romdata <= X"82006008";
    when 16#06C3# => romdata <= X"84102000";
    when 16#06C4# => romdata <= X"8528A003";
    when 16#06C5# => romdata <= X"03100031";
    when 16#06C6# => romdata <= X"8210636C";
    when 16#06C7# => romdata <= X"84004002";
    when 16#06C8# => romdata <= X"81C3E008";
    when 16#06C9# => romdata <= X"D000A004";
    when 16#06CA# => romdata <= X"9DE3BFA0";
    when 16#06CB# => romdata <= X"C2062084";
    when 16#06CC# => romdata <= X"C2006014";
    when 16#06CD# => romdata <= X"11100030";
    when 16#06CE# => romdata <= X"D20060FC";
    when 16#06CF# => romdata <= X"90122180";
    when 16#06D0# => romdata <= X"7FFFFE21";
    when 16#06D1# => romdata <= X"B0102000";
    when 16#06D2# => romdata <= X"81C7E008";
    when 16#06D3# => romdata <= X"81E80000";
    when 16#06D4# => romdata <= X"9DE3BFA0";
    when 16#06D5# => romdata <= X"11100030";
    when 16#06D6# => romdata <= X"7FFFFE1B";
    when 16#06D7# => romdata <= X"90122198";
    when 16#06D8# => romdata <= X"11100030";
    when 16#06D9# => romdata <= X"7FFFFE18";
    when 16#06DA# => romdata <= X"901221E0";
    when 16#06DB# => romdata <= X"11100030";
    when 16#06DC# => romdata <= X"7FFFFE15";
    when 16#06DD# => romdata <= X"90122208";
    when 16#06DE# => romdata <= X"11100030";
    when 16#06DF# => romdata <= X"7FFFFE12";
    when 16#06E0# => romdata <= X"90122220";
    when 16#06E1# => romdata <= X"11100030";
    when 16#06E2# => romdata <= X"7FFFFE0F";
    when 16#06E3# => romdata <= X"90122250";
    when 16#06E4# => romdata <= X"11100030";
    when 16#06E5# => romdata <= X"7FFFFE0C";
    when 16#06E6# => romdata <= X"90122278";
    when 16#06E7# => romdata <= X"11100030";
    when 16#06E8# => romdata <= X"7FFFFE09";
    when 16#06E9# => romdata <= X"901222A8";
    when 16#06EA# => romdata <= X"11100030";
    when 16#06EB# => romdata <= X"7FFFFE06";
    when 16#06EC# => romdata <= X"901222C0";
    when 16#06ED# => romdata <= X"11100030";
    when 16#06EE# => romdata <= X"7FFFFE03";
    when 16#06EF# => romdata <= X"901222F0";
    when 16#06F0# => romdata <= X"B2100018";
    when 16#06F1# => romdata <= X"31100030";
    when 16#06F2# => romdata <= X"7FFFFDFF";
    when 16#06F3# => romdata <= X"91EE2308";
    when 16#06F4# => romdata <= X"01000000";
    when 16#06F5# => romdata <= X"9DE3BFA0";
    when 16#06F6# => romdata <= X"11100030";
    when 16#06F7# => romdata <= X"7FFFFDFA";
    when 16#06F8# => romdata <= X"90122310";
    when 16#06F9# => romdata <= X"C2062084";
    when 16#06FA# => romdata <= X"25100030";
    when 16#06FB# => romdata <= X"A2102000";
    when 16#06FC# => romdata <= X"E0006018";
    when 16#06FD# => romdata <= X"A414A328";
    when 16#06FE# => romdata <= X"92100010";
    when 16#06FF# => romdata <= X"D4040000";
    when 16#0700# => romdata <= X"90100012";
    when 16#0701# => romdata <= X"7FFFFDF0";
    when 16#0702# => romdata <= X"A0042004";
    when 16#0703# => romdata <= X"7FFFFD68";
    when 16#0704# => romdata <= X"01000000";
    when 16#0705# => romdata <= X"80A22000";
    when 16#0706# => romdata <= X"12BFFFFD";
    when 16#0707# => romdata <= X"01000000";
    when 16#0708# => romdata <= X"A2046001";
    when 16#0709# => romdata <= X"80A46210";
    when 16#070A# => romdata <= X"12BFFFF5";
    when 16#070B# => romdata <= X"92100010";
    when 16#070C# => romdata <= X"81C7E008";
    when 16#070D# => romdata <= X"91E82000";
    when 16#070E# => romdata <= X"9DE3BFA0";
    when 16#070F# => romdata <= X"C2062084";
    when 16#0710# => romdata <= X"C2004000";
    when 16#0711# => romdata <= X"D2006FF0";
    when 16#0712# => romdata <= X"0300003F";
    when 16#0713# => romdata <= X"821063FF";
    when 16#0714# => romdata <= X"11100030";
    when 16#0715# => romdata <= X"920A4001";
    when 16#0716# => romdata <= X"7FFFFDDB";
    when 16#0717# => romdata <= X"90122338";
    when 16#0718# => romdata <= X"C2062084";
    when 16#0719# => romdata <= X"C2004000";
    when 16#071A# => romdata <= X"11100030";
    when 16#071B# => romdata <= X"D2106FF0";
    when 16#071C# => romdata <= X"90122360";
    when 16#071D# => romdata <= X"25100031";
    when 16#071E# => romdata <= X"2B100031";
    when 16#071F# => romdata <= X"A414A36C";
    when 16#0720# => romdata <= X"29100030";
    when 16#0721# => romdata <= X"27100030";
    when 16#0722# => romdata <= X"7FFFFDCF";
    when 16#0723# => romdata <= X"A0102000";
    when 16#0724# => romdata <= X"AA1563E4";
    when 16#0725# => romdata <= X"A8152378";
    when 16#0726# => romdata <= X"A614E388";
    when 16#0727# => romdata <= X"AC04A008";
    when 16#0728# => romdata <= X"C2062084";
    when 16#0729# => romdata <= X"C4004000";
    when 16#072A# => romdata <= X"832C2005";
    when 16#072B# => romdata <= X"C6008001";
    when 16#072C# => romdata <= X"80A0E000";
    when 16#072D# => romdata <= X"0280002A";
    when 16#072E# => romdata <= X"01000000";
    when 16#072F# => romdata <= X"DA008001";
    when 16#0730# => romdata <= X"C8008001";
    when 16#0731# => romdata <= X"E2008001";
    when 16#0732# => romdata <= X"8931200C";
    when 16#0733# => romdata <= X"88892FFF";
    when 16#0734# => romdata <= X"0280000C";
    when 16#0735# => romdata <= X"9B336018";
    when 16#0736# => romdata <= X"84100016";
    when 16#0737# => romdata <= X"82102001";
    when 16#0738# => romdata <= X"C6008000";
    when 16#0739# => romdata <= X"80A10003";
    when 16#073A# => romdata <= X"22800008";
    when 16#073B# => romdata <= X"83286003";
    when 16#073C# => romdata <= X"82006001";
    when 16#073D# => romdata <= X"80A0600F";
    when 16#073E# => romdata <= X"12BFFFFA";
    when 16#073F# => romdata <= X"8400A008";
    when 16#0740# => romdata <= X"82102000";
    when 16#0741# => romdata <= X"83286003";
    when 16#0742# => romdata <= X"80A36000";
    when 16#0743# => romdata <= X"82048001";
    when 16#0744# => romdata <= X"02800008";
    when 16#0745# => romdata <= X"D2006004";
    when 16#0746# => romdata <= X"80A36001";
    when 16#0747# => romdata <= X"02800006";
    when 16#0748# => romdata <= X"82102001";
    when 16#0749# => romdata <= X"80A360F1";
    when 16#074A# => romdata <= X"02800003";
    when 16#074B# => romdata <= X"82102002";
    when 16#074C# => romdata <= X"82102000";
    when 16#074D# => romdata <= X"83286003";
    when 16#074E# => romdata <= X"82054001";
    when 16#074F# => romdata <= X"90100014";
    when 16#0750# => romdata <= X"7FFFFDA1";
    when 16#0751# => romdata <= X"D4006004";
    when 16#0752# => romdata <= X"95346005";
    when 16#0753# => romdata <= X"90100013";
    when 16#0754# => romdata <= X"940AA01F";
    when 16#0755# => romdata <= X"7FFFFD9C";
    when 16#0756# => romdata <= X"92100010";
    when 16#0757# => romdata <= X"7FFFFD14";
    when 16#0758# => romdata <= X"01000000";
    when 16#0759# => romdata <= X"80A22000";
    when 16#075A# => romdata <= X"12BFFFFD";
    when 16#075B# => romdata <= X"01000000";
    when 16#075C# => romdata <= X"A0042001";
    when 16#075D# => romdata <= X"80A42010";
    when 16#075E# => romdata <= X"12BFFFCB";
    when 16#075F# => romdata <= X"C2062084";
    when 16#0760# => romdata <= X"2D100031";
    when 16#0761# => romdata <= X"39100031";
    when 16#0762# => romdata <= X"AC15A36C";
    when 16#0763# => romdata <= X"3B100030";
    when 16#0764# => romdata <= X"2F100030";
    when 16#0765# => romdata <= X"B81723E4";
    when 16#0766# => romdata <= X"BA176378";
    when 16#0767# => romdata <= X"AE15E3A8";
    when 16#0768# => romdata <= X"A2102000";
    when 16#0769# => romdata <= X"AA102000";
    when 16#076A# => romdata <= X"293FFC00";
    when 16#076B# => romdata <= X"B605A008";
    when 16#076C# => romdata <= X"84046040";
    when 16#076D# => romdata <= X"C2004000";
    when 16#076E# => romdata <= X"8528A005";
    when 16#076F# => romdata <= X"872C6005";
    when 16#0770# => romdata <= X"E4004002";
    when 16#0771# => romdata <= X"86004003";
    when 16#0772# => romdata <= X"E0004002";
    when 16#0773# => romdata <= X"E600E810";
    when 16#0774# => romdata <= X"F400E810";
    when 16#0775# => romdata <= X"C2004002";
    when 16#0776# => romdata <= X"A134200C";
    when 16#0777# => romdata <= X"80A06000";
    when 16#0778# => romdata <= X"A534A018";
    when 16#0779# => romdata <= X"A00C2FFF";
    when 16#077A# => romdata <= X"02800027";
    when 16#077B# => romdata <= X"A60CC014";
    when 16#077C# => romdata <= X"80A42000";
    when 16#077D# => romdata <= X"0280000B";
    when 16#077E# => romdata <= X"82102001";
    when 16#077F# => romdata <= X"8410001B";
    when 16#0780# => romdata <= X"C6008000";
    when 16#0781# => romdata <= X"80A40003";
    when 16#0782# => romdata <= X"22800008";
    when 16#0783# => romdata <= X"83286003";
    when 16#0784# => romdata <= X"82006001";
    when 16#0785# => romdata <= X"80A0600F";
    when 16#0786# => romdata <= X"12BFFFFA";
    when 16#0787# => romdata <= X"8400A008";
    when 16#0788# => romdata <= X"82102000";
    when 16#0789# => romdata <= X"83286003";
    when 16#078A# => romdata <= X"80A4A000";
    when 16#078B# => romdata <= X"82058001";
    when 16#078C# => romdata <= X"02800008";
    when 16#078D# => romdata <= X"D2006004";
    when 16#078E# => romdata <= X"80A4A001";
    when 16#078F# => romdata <= X"02800006";
    when 16#0790# => romdata <= X"82102001";
    when 16#0791# => romdata <= X"80A4A0F1";
    when 16#0792# => romdata <= X"02800003";
    when 16#0793# => romdata <= X"82102002";
    when 16#0794# => romdata <= X"82102000";
    when 16#0795# => romdata <= X"83286003";
    when 16#0796# => romdata <= X"82070001";
    when 16#0797# => romdata <= X"9010001D";
    when 16#0798# => romdata <= X"7FFFFD59";
    when 16#0799# => romdata <= X"D4006004";
    when 16#079A# => romdata <= X"B52EA010";
    when 16#079B# => romdata <= X"90100017";
    when 16#079C# => romdata <= X"960E8014";
    when 16#079D# => romdata <= X"92100011";
    when 16#079E# => romdata <= X"9634C00B";
    when 16#079F# => romdata <= X"7FFFFD52";
    when 16#07A0# => romdata <= X"94100013";
    when 16#07A1# => romdata <= X"80A42006";
    when 16#07A2# => romdata <= X"0280005B";
    when 16#07A3# => romdata <= X"80A4A001";
    when 16#07A4# => romdata <= X"7FFFFCC7";
    when 16#07A5# => romdata <= X"01000000";
    when 16#07A6# => romdata <= X"80A22000";
    when 16#07A7# => romdata <= X"12BFFFFD";
    when 16#07A8# => romdata <= X"01000000";
    when 16#07A9# => romdata <= X"A2046001";
    when 16#07AA# => romdata <= X"80A46010";
    when 16#07AB# => romdata <= X"32BFFFC1";
    when 16#07AC# => romdata <= X"C2062084";
    when 16#07AD# => romdata <= X"80A56000";
    when 16#07AE# => romdata <= X"0280004D";
    when 16#07AF# => romdata <= X"230003FF";
    when 16#07B0# => romdata <= X"25100031";
    when 16#07B1# => romdata <= X"AE1463FF";
    when 16#07B2# => romdata <= X"A414A36C";
    when 16#07B3# => romdata <= X"2D100031";
    when 16#07B4# => romdata <= X"29100030";
    when 16#07B5# => romdata <= X"27100030";
    when 16#07B6# => romdata <= X"AC15A3E4";
    when 16#07B7# => romdata <= X"A81523C8";
    when 16#07B8# => romdata <= X"A614E3D8";
    when 16#07B9# => romdata <= X"A0102000";
    when 16#07BA# => romdata <= X"A2146300";
    when 16#07BB# => romdata <= X"BA04A008";
    when 16#07BC# => romdata <= X"832C2003";
    when 16#07BD# => romdata <= X"C4062084";
    when 16#07BE# => romdata <= X"C400A004";
    when 16#07BF# => romdata <= X"D8008001";
    when 16#07C0# => romdata <= X"86008001";
    when 16#07C1# => romdata <= X"C8008001";
    when 16#07C2# => romdata <= X"DA00E004";
    when 16#07C3# => romdata <= X"F800E004";
    when 16#07C4# => romdata <= X"C2008001";
    when 16#07C5# => romdata <= X"80A06000";
    when 16#07C6# => romdata <= X"0280002C";
    when 16#07C7# => romdata <= X"8931200C";
    when 16#07C8# => romdata <= X"88892FFF";
    when 16#07C9# => romdata <= X"0280000B";
    when 16#07CA# => romdata <= X"8410001D";
    when 16#07CB# => romdata <= X"82102001";
    when 16#07CC# => romdata <= X"C6008000";
    when 16#07CD# => romdata <= X"80A10003";
    when 16#07CE# => romdata <= X"22800008";
    when 16#07CF# => romdata <= X"85332018";
    when 16#07D0# => romdata <= X"82006001";
    when 16#07D1# => romdata <= X"80A0600F";
    when 16#07D2# => romdata <= X"12BFFFFA";
    when 16#07D3# => romdata <= X"8400A008";
    when 16#07D4# => romdata <= X"82102000";
    when 16#07D5# => romdata <= X"85332018";
    when 16#07D6# => romdata <= X"83286003";
    when 16#07D7# => romdata <= X"80A0A000";
    when 16#07D8# => romdata <= X"82048001";
    when 16#07D9# => romdata <= X"02800008";
    when 16#07DA# => romdata <= X"D2006004";
    when 16#07DB# => romdata <= X"80A0A001";
    when 16#07DC# => romdata <= X"02800006";
    when 16#07DD# => romdata <= X"82102001";
    when 16#07DE# => romdata <= X"80A0A0F1";
    when 16#07DF# => romdata <= X"02800003";
    when 16#07E0# => romdata <= X"82102002";
    when 16#07E1# => romdata <= X"82102000";
    when 16#07E2# => romdata <= X"83286003";
    when 16#07E3# => romdata <= X"82058001";
    when 16#07E4# => romdata <= X"B7336010";
    when 16#07E5# => romdata <= X"D4006004";
    when 16#07E6# => romdata <= X"7FFFFD0B";
    when 16#07E7# => romdata <= X"90100014";
    when 16#07E8# => romdata <= X"B60EC011";
    when 16#07E9# => romdata <= X"972F2004";
    when 16#07EA# => romdata <= X"B615401B";
    when 16#07EB# => romdata <= X"960AC011";
    when 16#07EC# => romdata <= X"9410001B";
    when 16#07ED# => romdata <= X"962DC00B";
    when 16#07EE# => romdata <= X"90100013";
    when 16#07EF# => romdata <= X"9616C00B";
    when 16#07F0# => romdata <= X"7FFFFD01";
    when 16#07F1# => romdata <= X"92100010";
    when 16#07F2# => romdata <= X"7FFFFC79";
    when 16#07F3# => romdata <= X"01000000";
    when 16#07F4# => romdata <= X"80A22000";
    when 16#07F5# => romdata <= X"12BFFFFD";
    when 16#07F6# => romdata <= X"01000000";
    when 16#07F7# => romdata <= X"A0042001";
    when 16#07F8# => romdata <= X"80A42010";
    when 16#07F9# => romdata <= X"12BFFFC4";
    when 16#07FA# => romdata <= X"832C2003";
    when 16#07FB# => romdata <= X"81C7E008";
    when 16#07FC# => romdata <= X"91E82000";
    when 16#07FD# => romdata <= X"22BFFFA7";
    when 16#07FE# => romdata <= X"AA100013";
    when 16#07FF# => romdata <= X"30BFFFA5";
    when 16#0800# => romdata <= X"9DE3BFA0";
    when 16#0801# => romdata <= X"7FFFFD06";
    when 16#0802# => romdata <= X"23017D78";
    when 16#0803# => romdata <= X"11100030";
    when 16#0804# => romdata <= X"7FFFFCED";
    when 16#0805# => romdata <= X"901223F8";
    when 16#0806# => romdata <= X"C2062084";
    when 16#0807# => romdata <= X"C2006010";
    when 16#0808# => romdata <= X"A0102000";
    when 16#0809# => romdata <= X"C4006040";
    when 16#080A# => romdata <= X"A2146100";
    when 16#080B# => romdata <= X"8410A004";
    when 16#080C# => romdata <= X"C4206040";
    when 16#080D# => romdata <= X"7FFFFCF7";
    when 16#080E# => romdata <= X"01000000";
    when 16#080F# => romdata <= X"80A22009";
    when 16#0810# => romdata <= X"04800013";
    when 16#0811# => romdata <= X"80A40011";
    when 16#0812# => romdata <= X"C2062084";
    when 16#0813# => romdata <= X"C2006010";
    when 16#0814# => romdata <= X"C4006040";
    when 16#0815# => romdata <= X"8408BFFB";
    when 16#0816# => romdata <= X"C4206040";
    when 16#0817# => romdata <= X"7FFFFCED";
    when 16#0818# => romdata <= X"B0102000";
    when 16#0819# => romdata <= X"94100010";
    when 16#081A# => romdata <= X"92100008";
    when 16#081B# => romdata <= X"11100031";
    when 16#081C# => romdata <= X"7FFFFCD5";
    when 16#081D# => romdata <= X"90122018";
    when 16#081E# => romdata <= X"11100031";
    when 16#081F# => romdata <= X"7FFFFCD2";
    when 16#0820# => romdata <= X"90122038";
    when 16#0821# => romdata <= X"81C7E008";
    when 16#0822# => romdata <= X"81E80000";
    when 16#0823# => romdata <= X"22BFFFF0";
    when 16#0824# => romdata <= X"C2062084";
    when 16#0825# => romdata <= X"10BFFFE8";
    when 16#0826# => romdata <= X"A0042001";
    when 16#0827# => romdata <= X"9DE3BFA0";
    when 16#0828# => romdata <= X"7FFFFCDF";
    when 16#0829# => romdata <= X"01000000";
    when 16#082A# => romdata <= X"11100031";
    when 16#082B# => romdata <= X"7FFFFCC6";
    when 16#082C# => romdata <= X"90122058";
    when 16#082D# => romdata <= X"C2062084";
    when 16#082E# => romdata <= X"C2006010";
    when 16#082F# => romdata <= X"C4006040";
    when 16#0830# => romdata <= X"8410A010";
    when 16#0831# => romdata <= X"23017D78";
    when 16#0832# => romdata <= X"C4206040";
    when 16#0833# => romdata <= X"7FFFFCD1";
    when 16#0834# => romdata <= X"A0102000";
    when 16#0835# => romdata <= X"80A22009";
    when 16#0836# => romdata <= X"1480000A";
    when 16#0837# => romdata <= X"A2146100";
    when 16#0838# => romdata <= X"80A40011";
    when 16#0839# => romdata <= X"22800008";
    when 16#083A# => romdata <= X"C2062084";
    when 16#083B# => romdata <= X"7FFFFCC9";
    when 16#083C# => romdata <= X"A0042001";
    when 16#083D# => romdata <= X"80A22009";
    when 16#083E# => romdata <= X"04BFFFFB";
    when 16#083F# => romdata <= X"80A40011";
    when 16#0840# => romdata <= X"C2062084";
    when 16#0841# => romdata <= X"C2006010";
    when 16#0842# => romdata <= X"C4006040";
    when 16#0843# => romdata <= X"8408BFEF";
    when 16#0844# => romdata <= X"C4206040";
    when 16#0845# => romdata <= X"7FFFFCBF";
    when 16#0846# => romdata <= X"B0102000";
    when 16#0847# => romdata <= X"92100008";
    when 16#0848# => romdata <= X"11100031";
    when 16#0849# => romdata <= X"7FFFFCA8";
    when 16#084A# => romdata <= X"90122078";
    when 16#084B# => romdata <= X"11100031";
    when 16#084C# => romdata <= X"7FFFFCA5";
    when 16#084D# => romdata <= X"90122098";
    when 16#084E# => romdata <= X"81C7E008";
    when 16#084F# => romdata <= X"81E80000";
    when 16#0850# => romdata <= X"9DE3BFA0";
    when 16#0851# => romdata <= X"13100031";
    when 16#0852# => romdata <= X"90100019";
    when 16#0853# => romdata <= X"921260B8";
    when 16#0854# => romdata <= X"40000119";
    when 16#0855# => romdata <= X"A0102000";
    when 16#0856# => romdata <= X"80A22000";
    when 16#0857# => romdata <= X"12800005";
    when 16#0858# => romdata <= X"90100019";
    when 16#0859# => romdata <= X"82102001";
    when 16#085A# => romdata <= X"A0102001";
    when 16#085B# => romdata <= X"C2262080";
    when 16#085C# => romdata <= X"13100031";
    when 16#085D# => romdata <= X"40000110";
    when 16#085E# => romdata <= X"921260C0";
    when 16#085F# => romdata <= X"80A22000";
    when 16#0860# => romdata <= X"12800005";
    when 16#0861# => romdata <= X"90100019";
    when 16#0862# => romdata <= X"82102002";
    when 16#0863# => romdata <= X"A0102002";
    when 16#0864# => romdata <= X"C2262080";
    when 16#0865# => romdata <= X"13100031";
    when 16#0866# => romdata <= X"40000107";
    when 16#0867# => romdata <= X"921260C8";
    when 16#0868# => romdata <= X"80A22000";
    when 16#0869# => romdata <= X"12800005";
    when 16#086A# => romdata <= X"90100019";
    when 16#086B# => romdata <= X"82102003";
    when 16#086C# => romdata <= X"A0102003";
    when 16#086D# => romdata <= X"C2262080";
    when 16#086E# => romdata <= X"13100031";
    when 16#086F# => romdata <= X"400000FE";
    when 16#0870# => romdata <= X"921260D0";
    when 16#0871# => romdata <= X"80A22000";
    when 16#0872# => romdata <= X"12800005";
    when 16#0873# => romdata <= X"90100019";
    when 16#0874# => romdata <= X"82102004";
    when 16#0875# => romdata <= X"A0102004";
    when 16#0876# => romdata <= X"C2262080";
    when 16#0877# => romdata <= X"13100031";
    when 16#0878# => romdata <= X"400000F5";
    when 16#0879# => romdata <= X"921260D8";
    when 16#087A# => romdata <= X"80A22000";
    when 16#087B# => romdata <= X"12800005";
    when 16#087C# => romdata <= X"90100019";
    when 16#087D# => romdata <= X"82102005";
    when 16#087E# => romdata <= X"A0102005";
    when 16#087F# => romdata <= X"C2262080";
    when 16#0880# => romdata <= X"13100031";
    when 16#0881# => romdata <= X"400000EC";
    when 16#0882# => romdata <= X"921260E0";
    when 16#0883# => romdata <= X"80A22000";
    when 16#0884# => romdata <= X"12800005";
    when 16#0885# => romdata <= X"90100019";
    when 16#0886# => romdata <= X"82102006";
    when 16#0887# => romdata <= X"A0102006";
    when 16#0888# => romdata <= X"C2262080";
    when 16#0889# => romdata <= X"13100031";
    when 16#088A# => romdata <= X"400000E3";
    when 16#088B# => romdata <= X"921260E8";
    when 16#088C# => romdata <= X"80A22000";
    when 16#088D# => romdata <= X"12800004";
    when 16#088E# => romdata <= X"82102007";
    when 16#088F# => romdata <= X"A0102007";
    when 16#0890# => romdata <= X"C2262080";
    when 16#0891# => romdata <= X"81C7E008";
    when 16#0892# => romdata <= X"91E80010";
    when 16#0893# => romdata <= X"9DE3BFA0";
    when 16#0894# => romdata <= X"25100006";
    when 16#0895# => romdata <= X"27100030";
    when 16#0896# => romdata <= X"29100031";
    when 16#0897# => romdata <= X"23100031";
    when 16#0898# => romdata <= X"A414A274";
    when 16#0899# => romdata <= X"A614E180";
    when 16#089A# => romdata <= X"A81520F0";
    when 16#089B# => romdata <= X"A2146108";
    when 16#089C# => romdata <= X"C20E0000";
    when 16#089D# => romdata <= X"83286018";
    when 16#089E# => romdata <= X"83386018";
    when 16#089F# => romdata <= X"80A06072";
    when 16#08A0# => romdata <= X"0280000B";
    when 16#08A1# => romdata <= X"80A42007";
    when 16#08A2# => romdata <= X"7FFFFE32";
    when 16#08A3# => romdata <= X"90100018";
    when 16#08A4# => romdata <= X"7FFFFC32";
    when 16#08A5# => romdata <= X"90100018";
    when 16#08A6# => romdata <= X"90100018";
    when 16#08A7# => romdata <= X"7FFFFFA9";
    when 16#08A8# => romdata <= X"92100018";
    when 16#08A9# => romdata <= X"A0100008";
    when 16#08AA# => romdata <= X"80A42007";
    when 16#08AB# => romdata <= X"0880000F";
    when 16#08AC# => romdata <= X"832C2002";
    when 16#08AD# => romdata <= X"90100014";
    when 16#08AE# => romdata <= X"7FFFFC43";
    when 16#08AF# => romdata <= X"92100018";
    when 16#08B0# => romdata <= X"82102000";
    when 16#08B1# => romdata <= X"83286018";
    when 16#08B2# => romdata <= X"83386018";
    when 16#08B3# => romdata <= X"80A06072";
    when 16#08B4# => romdata <= X"12BFFFEE";
    when 16#08B5# => romdata <= X"C02E0000";
    when 16#08B6# => romdata <= X"80A42007";
    when 16#08B7# => romdata <= X"18BFFFF7";
    when 16#08B8# => romdata <= X"90100014";
    when 16#08B9# => romdata <= X"832C2002";
    when 16#08BA# => romdata <= X"C2048001";
    when 16#08BB# => romdata <= X"81C04000";
    when 16#08BC# => romdata <= X"01000000";
    when 16#08BD# => romdata <= X"C2062084";
    when 16#08BE# => romdata <= X"C2006014";
    when 16#08BF# => romdata <= X"90100013";
    when 16#08C0# => romdata <= X"D20060FC";
    when 16#08C1# => romdata <= X"7FFFFC30";
    when 16#08C2# => romdata <= X"A0102007";
    when 16#08C3# => romdata <= X"7FFFFE4B";
    when 16#08C4# => romdata <= X"90100018";
    when 16#08C5# => romdata <= X"7FFFFF62";
    when 16#08C6# => romdata <= X"90100018";
    when 16#08C7# => romdata <= X"7FFFFF39";
    when 16#08C8# => romdata <= X"90100018";
    when 16#08C9# => romdata <= X"7FFFFE2C";
    when 16#08CA# => romdata <= X"90100018";
    when 16#08CB# => romdata <= X"7FFFFD2E";
    when 16#08CC# => romdata <= X"90100018";
    when 16#08CD# => romdata <= X"7FFFFC24";
    when 16#08CE# => romdata <= X"90100011";
    when 16#08CF# => romdata <= X"7FFFFC07";
    when 16#08D0# => romdata <= X"90100018";
    when 16#08D1# => romdata <= X"10BFFFCC";
    when 16#08D2# => romdata <= X"C20E0000";
    when 16#08D3# => romdata <= X"7FFFFE22";
    when 16#08D4# => romdata <= X"90100018";
    when 16#08D5# => romdata <= X"30BFFFF8";
    when 16#08D6# => romdata <= X"7FFFFF2A";
    when 16#08D7# => romdata <= X"90100018";
    when 16#08D8# => romdata <= X"30BFFFF5";
    when 16#08D9# => romdata <= X"7FFFFF4E";
    when 16#08DA# => romdata <= X"90100018";
    when 16#08DB# => romdata <= X"30BFFFF2";
    when 16#08DC# => romdata <= X"7FFFFE32";
    when 16#08DD# => romdata <= X"90100018";
    when 16#08DE# => romdata <= X"30BFFFEF";
    when 16#08DF# => romdata <= X"C2062084";
    when 16#08E0# => romdata <= X"C2006014";
    when 16#08E1# => romdata <= X"90100013";
    when 16#08E2# => romdata <= X"D20060FC";
    when 16#08E3# => romdata <= X"7FFFFC0E";
    when 16#08E4# => romdata <= X"01000000";
    when 16#08E5# => romdata <= X"30BFFFE8";
    when 16#08E6# => romdata <= X"81C3E008";
    when 16#08E7# => romdata <= X"01000000";
    when 16#08E8# => romdata <= X"81C3E008";
    when 16#08E9# => romdata <= X"01000000";
    when 16#08EA# => romdata <= X"81C3E008";
    when 16#08EB# => romdata <= X"01000000";
    when 16#08EC# => romdata <= X"81C3E008";
    when 16#08ED# => romdata <= X"01000000";
    when 16#08EE# => romdata <= X"03200000";
    when 16#08EF# => romdata <= X"84106200";
    when 16#08F0# => romdata <= X"C4222010";
    when 16#08F1# => romdata <= X"84103000";
    when 16#08F2# => romdata <= X"C4220000";
    when 16#08F3# => romdata <= X"052003FC";
    when 16#08F4# => romdata <= X"C4222004";
    when 16#08F5# => romdata <= X"84106100";
    when 16#08F6# => romdata <= X"82106300";
    when 16#08F7# => romdata <= X"C222200C";
    when 16#08F8# => romdata <= X"03200001";
    when 16#08F9# => romdata <= X"C4222008";
    when 16#08FA# => romdata <= X"C2222014";
    when 16#08FB# => romdata <= X"03340000";
    when 16#08FC# => romdata <= X"81C3E008";
    when 16#08FD# => romdata <= X"C2222018";
    when 16#08FE# => romdata <= X"11100008";
    when 16#08FF# => romdata <= X"13100037";
    when 16#0900# => romdata <= X"15100032";
    when 16#0901# => romdata <= X"901223B0";
    when 16#0902# => romdata <= X"921261B8";
    when 16#0903# => romdata <= X"9412A2BC";
    when 16#0904# => romdata <= X"8213C000";
    when 16#0905# => romdata <= X"4000005F";
    when 16#0906# => romdata <= X"9E104000";
    when 16#0907# => romdata <= X"01000000";
    when 16#0908# => romdata <= X"9DE3BFA0";
    when 16#0909# => romdata <= X"84102047";
    when 16#090A# => romdata <= X"C2062008";
    when 16#090B# => romdata <= X"C420600C";
    when 16#090C# => romdata <= X"05000010";
    when 16#090D# => romdata <= X"8410A003";
    when 16#090E# => romdata <= X"C4206008";
    when 16#090F# => romdata <= X"C206200C";
    when 16#0910# => romdata <= X"84102042";
    when 16#0911# => romdata <= X"C4206004";
    when 16#0912# => romdata <= X"C4204000";
    when 16#0913# => romdata <= X"C0206018";
    when 16#0914# => romdata <= X"C0206028";
    when 16#0915# => romdata <= X"050003D0";
    when 16#0916# => romdata <= X"8410A240";
    when 16#0917# => romdata <= X"C4206014";
    when 16#0918# => romdata <= X"8410200F";
    when 16#0919# => romdata <= X"C4206018";
    when 16#091A# => romdata <= X"0300FBC5";
    when 16#091B# => romdata <= X"82106080";
    when 16#091C# => romdata <= X"C8062018";
    when 16#091D# => romdata <= X"84102000";
    when 16#091E# => romdata <= X"C2212800";
    when 16#091F# => romdata <= X"1B3FC48D";
    when 16#0920# => romdata <= X"82102000";
    when 16#0921# => romdata <= X"8400800D";
    when 16#0922# => romdata <= X"87286006";
    when 16#0923# => romdata <= X"C4210003";
    when 16#0924# => romdata <= X"82006001";
    when 16#0925# => romdata <= X"80A06020";
    when 16#0926# => romdata <= X"12BFFFFB";
    when 16#0927# => romdata <= X"84100001";
    when 16#0928# => romdata <= X"C2062010";
    when 16#0929# => romdata <= X"C0204000";
    when 16#092A# => romdata <= X"C0206040";
    when 16#092B# => romdata <= X"84103FFF";
    when 16#092C# => romdata <= X"92102004";
    when 16#092D# => romdata <= X"C420600C";
    when 16#092E# => romdata <= X"11100005";
    when 16#092F# => romdata <= X"4000209A";
    when 16#0930# => romdata <= X"90122064";
    when 16#0931# => romdata <= X"92102003";
    when 16#0932# => romdata <= X"11100005";
    when 16#0933# => romdata <= X"40002096";
    when 16#0934# => romdata <= X"90122028";
    when 16#0935# => romdata <= X"92102002";
    when 16#0936# => romdata <= X"11100005";
    when 16#0937# => romdata <= X"40002092";
    when 16#0938# => romdata <= X"90122038";
    when 16#0939# => romdata <= X"C2062010";
    when 16#093A# => romdata <= X"C4006040";
    when 16#093B# => romdata <= X"8410A008";
    when 16#093C# => romdata <= X"C4206040";
    when 16#093D# => romdata <= X"81C7E008";
    when 16#093E# => romdata <= X"81E80000";
    when 16#093F# => romdata <= X"9DE3BFA0";
    when 16#0940# => romdata <= X"33100037";
    when 16#0941# => romdata <= X"9016625C";
    when 16#0942# => romdata <= X"31100008";
    when 16#0943# => romdata <= X"B2100008";
    when 16#0944# => romdata <= X"7FFFFFA4";
    when 16#0945# => romdata <= X"35100032";
    when 16#0946# => romdata <= X"B01623B0";
    when 16#0947# => romdata <= X"4000001D";
    when 16#0948# => romdata <= X"95EEA2BC";
    when 16#0949# => romdata <= X"01000000";
    when 16#094A# => romdata <= X"9DE3BFA0";
    when 16#094B# => romdata <= X"21100037";
    when 16#094C# => romdata <= X"7FFFFFA2";
    when 16#094D# => romdata <= X"9014225C";
    when 16#094E# => romdata <= X"7FFFFFBA";
    when 16#094F# => romdata <= X"9014225C";
    when 16#0950# => romdata <= X"A014225C";
    when 16#0951# => romdata <= X"7FFFFB17";
    when 16#0952# => romdata <= X"D0042008";
    when 16#0953# => romdata <= X"92100010";
    when 16#0954# => romdata <= X"21100037";
    when 16#0955# => romdata <= X"7FFFFD50";
    when 16#0956# => romdata <= X"901421D4";
    when 16#0957# => romdata <= X"901421D4";
    when 16#0958# => romdata <= X"7FFFFF3B";
    when 16#0959# => romdata <= X"B0102000";
    when 16#095A# => romdata <= X"81C7E008";
    when 16#095B# => romdata <= X"81E80000";
    when 16#095C# => romdata <= X"92100008";
    when 16#095D# => romdata <= X"94102000";
    when 16#095E# => romdata <= X"90102000";
    when 16#095F# => romdata <= X"96102000";
    when 16#0960# => romdata <= X"8213C000";
    when 16#0961# => romdata <= X"4000006F";
    when 16#0962# => romdata <= X"9E104000";
    when 16#0963# => romdata <= X"01000000";
    when 16#0964# => romdata <= X"82100009";
    when 16#0965# => romdata <= X"9610000A";
    when 16#0966# => romdata <= X"92100008";
    when 16#0967# => romdata <= X"94100001";
    when 16#0968# => romdata <= X"90102002";
    when 16#0969# => romdata <= X"8213C000";
    when 16#096A# => romdata <= X"40000066";
    when 16#096B# => romdata <= X"9E104000";
    when 16#096C# => romdata <= X"01000000";
    when 16#096D# => romdata <= X"82124008";
    when 16#096E# => romdata <= X"80886003";
    when 16#096F# => romdata <= X"3280001E";
    when 16#0970# => romdata <= X"C24A0000";
    when 16#0971# => romdata <= X"C2020000";
    when 16#0972# => romdata <= X"C4024000";
    when 16#0973# => romdata <= X"80A04002";
    when 16#0974# => romdata <= X"12800018";
    when 16#0975# => romdata <= X"053FBFBF";
    when 16#0976# => romdata <= X"07202020";
    when 16#0977# => romdata <= X"8410A2FF";
    when 16#0978# => romdata <= X"8610E080";
    when 16#0979# => romdata <= X"88100002";
    when 16#097A# => romdata <= X"84004002";
    when 16#097B# => romdata <= X"82288001";
    when 16#097C# => romdata <= X"80884003";
    when 16#097D# => romdata <= X"22800009";
    when 16#097E# => romdata <= X"90022004";
    when 16#097F# => romdata <= X"81C3E008";
    when 16#0980# => romdata <= X"90102000";
    when 16#0981# => romdata <= X"82288001";
    when 16#0982# => romdata <= X"80884003";
    when 16#0983# => romdata <= X"32800022";
    when 16#0984# => romdata <= X"90102000";
    when 16#0985# => romdata <= X"90022004";
    when 16#0986# => romdata <= X"92026004";
    when 16#0987# => romdata <= X"C2020000";
    when 16#0988# => romdata <= X"C4024000";
    when 16#0989# => romdata <= X"80A04002";
    when 16#098A# => romdata <= X"02BFFFF7";
    when 16#098B# => romdata <= X"84004004";
    when 16#098C# => romdata <= X"C24A0000";
    when 16#098D# => romdata <= X"80A06000";
    when 16#098E# => romdata <= X"1280000A";
    when 16#098F# => romdata <= X"C60A0000";
    when 16#0990# => romdata <= X"10800011";
    when 16#0991# => romdata <= X"C20A4000";
    when 16#0992# => romdata <= X"90022001";
    when 16#0993# => romdata <= X"C24A0000";
    when 16#0994# => romdata <= X"92026001";
    when 16#0995# => romdata <= X"80A06000";
    when 16#0996# => romdata <= X"0280000A";
    when 16#0997# => romdata <= X"C60A0000";
    when 16#0998# => romdata <= X"C44A4000";
    when 16#0999# => romdata <= X"80A04002";
    when 16#099A# => romdata <= X"02BFFFF8";
    when 16#099B# => romdata <= X"C20A4000";
    when 16#099C# => romdata <= X"8608E0FF";
    when 16#099D# => romdata <= X"820860FF";
    when 16#099E# => romdata <= X"81C3E008";
    when 16#099F# => romdata <= X"9020C001";
    when 16#09A0# => romdata <= X"C20A4000";
    when 16#09A1# => romdata <= X"8608E0FF";
    when 16#09A2# => romdata <= X"820860FF";
    when 16#09A3# => romdata <= X"81C3E008";
    when 16#09A4# => romdata <= X"9020C001";
    when 16#09A5# => romdata <= X"81C3E008";
    when 16#09A6# => romdata <= X"01000000";
    when 16#09A7# => romdata <= X"9DE3BED0";
    when 16#09A8# => romdata <= X"82102208";
    when 16#09A9# => romdata <= X"C237BF40";
    when 16#09AA# => romdata <= X"031FFFFF";
    when 16#09AB# => romdata <= X"821063FF";
    when 16#09AC# => romdata <= X"C227BF48";
    when 16#09AD# => romdata <= X"C227BF3C";
    when 16#09AE# => romdata <= X"82103FFF";
    when 16#09AF# => romdata <= X"F227BF44";
    when 16#09B0# => romdata <= X"C237BF42";
    when 16#09B1# => romdata <= X"90100018";
    when 16#09B2# => romdata <= X"F227BF34";
    when 16#09B3# => romdata <= X"9410001A";
    when 16#09B4# => romdata <= X"9610001B";
    when 16#09B5# => romdata <= X"400002AD";
    when 16#09B6# => romdata <= X"9207BF34";
    when 16#09B7# => romdata <= X"C207BF34";
    when 16#09B8# => romdata <= X"C0284000";
    when 16#09B9# => romdata <= X"81C7E008";
    when 16#09BA# => romdata <= X"91E80008";
    when 16#09BB# => romdata <= X"9DE3BED0";
    when 16#09BC# => romdata <= X"03100032";
    when 16#09BD# => romdata <= X"D00062C8";
    when 16#09BE# => romdata <= X"82102208";
    when 16#09BF# => romdata <= X"C237BF40";
    when 16#09C0# => romdata <= X"031FFFFF";
    when 16#09C1# => romdata <= X"821063FF";
    when 16#09C2# => romdata <= X"C227BF48";
    when 16#09C3# => romdata <= X"C227BF3C";
    when 16#09C4# => romdata <= X"82103FFF";
    when 16#09C5# => romdata <= X"F027BF44";
    when 16#09C6# => romdata <= X"F027BF34";
    when 16#09C7# => romdata <= X"C237BF42";
    when 16#09C8# => romdata <= X"94100019";
    when 16#09C9# => romdata <= X"9610001A";
    when 16#09CA# => romdata <= X"40000298";
    when 16#09CB# => romdata <= X"9207BF34";
    when 16#09CC# => romdata <= X"C207BF34";
    when 16#09CD# => romdata <= X"C0284000";
    when 16#09CE# => romdata <= X"81C7E008";
    when 16#09CF# => romdata <= X"91E80008";
    when 16#09D0# => romdata <= X"9DE3BFA0";
    when 16#09D1# => romdata <= X"21100037";
    when 16#09D2# => romdata <= X"400020D2";
    when 16#09D3# => romdata <= X"9014227C";
    when 16#09D4# => romdata <= X"03100031";
    when 16#09D5# => romdata <= X"E20063FC";
    when 16#09D6# => romdata <= X"D0046148";
    when 16#09D7# => romdata <= X"80A22000";
    when 16#09D8# => romdata <= X"2280003D";
    when 16#09D9# => romdata <= X"9004614C";
    when 16#09DA# => romdata <= X"C2022004";
    when 16#09DB# => romdata <= X"80A0601F";
    when 16#09DC# => romdata <= X"1480001E";
    when 16#09DD# => romdata <= X"01000000";
    when 16#09DE# => romdata <= X"80A62000";
    when 16#09DF# => romdata <= X"02800012";
    when 16#09E0# => romdata <= X"84006002";
    when 16#09E1# => romdata <= X"C4022004";
    when 16#09E2# => romdata <= X"82006022";
    when 16#09E3# => romdata <= X"8600A042";
    when 16#09E4# => romdata <= X"89286002";
    when 16#09E5# => romdata <= X"8728E002";
    when 16#09E6# => romdata <= X"C2022188";
    when 16#09E7# => romdata <= X"F4220004";
    when 16#09E8# => romdata <= X"F6220003";
    when 16#09E9# => romdata <= X"86102001";
    when 16#09EA# => romdata <= X"8728C002";
    when 16#09EB# => romdata <= X"82104003";
    when 16#09EC# => romdata <= X"C2222188";
    when 16#09ED# => romdata <= X"80A62002";
    when 16#09EE# => romdata <= X"02800019";
    when 16#09EF# => romdata <= X"82100002";
    when 16#09F0# => romdata <= X"84006002";
    when 16#09F1# => romdata <= X"8528A002";
    when 16#09F2# => romdata <= X"82006001";
    when 16#09F3# => romdata <= X"C2222004";
    when 16#09F4# => romdata <= X"F2220002";
    when 16#09F5# => romdata <= X"B0102000";
    when 16#09F6# => romdata <= X"400020C4";
    when 16#09F7# => romdata <= X"9014227C";
    when 16#09F8# => romdata <= X"81C7E008";
    when 16#09F9# => romdata <= X"81E80000";
    when 16#09FA# => romdata <= X"40000028";
    when 16#09FB# => romdata <= X"90102190";
    when 16#09FC# => romdata <= X"80A22000";
    when 16#09FD# => romdata <= X"2280001A";
    when 16#09FE# => romdata <= X"9014227C";
    when 16#09FF# => romdata <= X"C2046148";
    when 16#0A00# => romdata <= X"C2220000";
    when 16#0A01# => romdata <= X"D0246148";
    when 16#0A02# => romdata <= X"C0222004";
    when 16#0A03# => romdata <= X"C0222188";
    when 16#0A04# => romdata <= X"C022218C";
    when 16#0A05# => romdata <= X"10BFFFD9";
    when 16#0A06# => romdata <= X"82102000";
    when 16#0A07# => romdata <= X"C202218C";
    when 16#0A08# => romdata <= X"86104003";
    when 16#0A09# => romdata <= X"82100002";
    when 16#0A0A# => romdata <= X"84006002";
    when 16#0A0B# => romdata <= X"8528A002";
    when 16#0A0C# => romdata <= X"C622218C";
    when 16#0A0D# => romdata <= X"82006001";
    when 16#0A0E# => romdata <= X"F2220002";
    when 16#0A0F# => romdata <= X"C2222004";
    when 16#0A10# => romdata <= X"B0102000";
    when 16#0A11# => romdata <= X"400020A9";
    when 16#0A12# => romdata <= X"9014227C";
    when 16#0A13# => romdata <= X"81C7E008";
    when 16#0A14# => romdata <= X"81E80000";
    when 16#0A15# => romdata <= X"10BFFFC5";
    when 16#0A16# => romdata <= X"D0246148";
    when 16#0A17# => romdata <= X"400020A3";
    when 16#0A18# => romdata <= X"B0103FFF";
    when 16#0A19# => romdata <= X"81C7E008";
    when 16#0A1A# => romdata <= X"81E80000";
    when 16#0A1B# => romdata <= X"92100008";
    when 16#0A1C# => romdata <= X"03100032";
    when 16#0A1D# => romdata <= X"D00062C8";
    when 16#0A1E# => romdata <= X"8213C000";
    when 16#0A1F# => romdata <= X"40001218";
    when 16#0A20# => romdata <= X"9E104000";
    when 16#0A21# => romdata <= X"01000000";
    when 16#0A22# => romdata <= X"92100008";
    when 16#0A23# => romdata <= X"03100032";
    when 16#0A24# => romdata <= X"D00062C8";
    when 16#0A25# => romdata <= X"8213C000";
    when 16#0A26# => romdata <= X"40000003";
    when 16#0A27# => romdata <= X"9E104000";
    when 16#0A28# => romdata <= X"01000000";
    when 16#0A29# => romdata <= X"9DE3BFA0";
    when 16#0A2A# => romdata <= X"84102000";
    when 16#0A2B# => romdata <= X"8206600B";
    when 16#0A2C# => romdata <= X"80A06016";
    when 16#0A2D# => romdata <= X"08800004";
    when 16#0A2E# => romdata <= X"A0102010";
    when 16#0A2F# => romdata <= X"A0087FF8";
    when 16#0A30# => romdata <= X"8534201F";
    when 16#0A31# => romdata <= X"80A40019";
    when 16#0A32# => romdata <= X"0A800046";
    when 16#0A33# => romdata <= X"8088A0FF";
    when 16#0A34# => romdata <= X"12800044";
    when 16#0A35# => romdata <= X"01000000";
    when 16#0A36# => romdata <= X"400001AF";
    when 16#0A37# => romdata <= X"90100018";
    when 16#0A38# => romdata <= X"80A421F7";
    when 16#0A39# => romdata <= X"18800041";
    when 16#0A3A# => romdata <= X"83342009";
    when 16#0A3B# => romdata <= X"23100034";
    when 16#0A3C# => romdata <= X"A2146020";
    when 16#0A3D# => romdata <= X"82044010";
    when 16#0A3E# => romdata <= X"E400600C";
    when 16#0A3F# => romdata <= X"80A48001";
    when 16#0A40# => romdata <= X"0280010F";
    when 16#0A41# => romdata <= X"99342003";
    when 16#0A42# => romdata <= X"C604A004";
    when 16#0A43# => romdata <= X"C404A00C";
    when 16#0A44# => romdata <= X"C204A008";
    when 16#0A45# => romdata <= X"8608FFFC";
    when 16#0A46# => romdata <= X"86048003";
    when 16#0A47# => romdata <= X"C800E004";
    when 16#0A48# => romdata <= X"88112001";
    when 16#0A49# => romdata <= X"C220A008";
    when 16#0A4A# => romdata <= X"C820E004";
    when 16#0A4B# => romdata <= X"C420600C";
    when 16#0A4C# => romdata <= X"90100018";
    when 16#0A4D# => romdata <= X"40000192";
    when 16#0A4E# => romdata <= X"B004A008";
    when 16#0A4F# => romdata <= X"81C7E008";
    when 16#0A50# => romdata <= X"81E80000";
    when 16#0A51# => romdata <= X"E6046008";
    when 16#0A52# => romdata <= X"E804E004";
    when 16#0A53# => romdata <= X"A80D3FFC";
    when 16#0A54# => romdata <= X"82250010";
    when 16#0A55# => romdata <= X"80A0600F";
    when 16#0A56# => romdata <= X"148000D2";
    when 16#0A57# => romdata <= X"80A40014";
    when 16#0A58# => romdata <= X"03100037";
    when 16#0A59# => romdata <= X"2F100035";
    when 16#0A5A# => romdata <= X"EA0062F0";
    when 16#0A5B# => romdata <= X"C205E02C";
    when 16#0A5C# => romdata <= X"AA056010";
    when 16#0A5D# => romdata <= X"80A07FFF";
    when 16#0A5E# => romdata <= X"02800004";
    when 16#0A5F# => romdata <= X"AA054010";
    when 16#0A60# => romdata <= X"AA056FFF";
    when 16#0A61# => romdata <= X"AA0D7000";
    when 16#0A62# => romdata <= X"90100018";
    when 16#0A63# => romdata <= X"40000188";
    when 16#0A64# => romdata <= X"92100015";
    when 16#0A65# => romdata <= X"80A23FFF";
    when 16#0A66# => romdata <= X"02800009";
    when 16#0A67# => romdata <= X"A4100008";
    when 16#0A68# => romdata <= X"8404C014";
    when 16#0A69# => romdata <= X"80A08008";
    when 16#0A6A# => romdata <= X"088000EC";
    when 16#0A6B# => romdata <= X"2D100037";
    when 16#0A6C# => romdata <= X"80A44013";
    when 16#0A6D# => romdata <= X"028000EA";
    when 16#0A6E# => romdata <= X"C205A2FC";
    when 16#0A6F# => romdata <= X"C2046008";
    when 16#0A70# => romdata <= X"C4006004";
    when 16#0A71# => romdata <= X"8408BFFC";
    when 16#0A72# => romdata <= X"82208010";
    when 16#0A73# => romdata <= X"80A0600F";
    when 16#0A74# => romdata <= X"14800122";
    when 16#0A75# => romdata <= X"80A40002";
    when 16#0A76# => romdata <= X"40000169";
    when 16#0A77# => romdata <= X"90100018";
    when 16#0A78# => romdata <= X"81C7E008";
    when 16#0A79# => romdata <= X"91E82000";
    when 16#0A7A# => romdata <= X"99342003";
    when 16#0A7B# => romdata <= X"80A06000";
    when 16#0A7C# => romdata <= X"0280000F";
    when 16#0A7D# => romdata <= X"872B2003";
    when 16#0A7E# => romdata <= X"80A06004";
    when 16#0A7F# => romdata <= X"08800092";
    when 16#0A80# => romdata <= X"99342006";
    when 16#0A81# => romdata <= X"9800605B";
    when 16#0A82# => romdata <= X"80A06014";
    when 16#0A83# => romdata <= X"08800008";
    when 16#0A84# => romdata <= X"872B2003";
    when 16#0A85# => romdata <= X"80A06054";
    when 16#0A86# => romdata <= X"18800113";
    when 16#0A87# => romdata <= X"80A06154";
    when 16#0A88# => romdata <= X"9934200C";
    when 16#0A89# => romdata <= X"9803206E";
    when 16#0A8A# => romdata <= X"872B2003";
    when 16#0A8B# => romdata <= X"23100034";
    when 16#0A8C# => romdata <= X"A2146020";
    when 16#0A8D# => romdata <= X"86044003";
    when 16#0A8E# => romdata <= X"E400E00C";
    when 16#0A8F# => romdata <= X"80A0C012";
    when 16#0A90# => romdata <= X"3280000B";
    when 16#0A91# => romdata <= X"C404A004";
    when 16#0A92# => romdata <= X"10800010";
    when 16#0A93# => romdata <= X"98032001";
    when 16#0A94# => romdata <= X"36800068";
    when 16#0A95# => romdata <= X"C604A00C";
    when 16#0A96# => romdata <= X"E404A00C";
    when 16#0A97# => romdata <= X"80A0C012";
    when 16#0A98# => romdata <= X"2280000A";
    when 16#0A99# => romdata <= X"98032001";
    when 16#0A9A# => romdata <= X"C404A004";
    when 16#0A9B# => romdata <= X"8408BFFC";
    when 16#0A9C# => romdata <= X"82208010";
    when 16#0A9D# => romdata <= X"80A0600F";
    when 16#0A9E# => romdata <= X"04BFFFF6";
    when 16#0A9F# => romdata <= X"80A06000";
    when 16#0AA0# => romdata <= X"98033FFF";
    when 16#0AA1# => romdata <= X"98032001";
    when 16#0AA2# => romdata <= X"07100034";
    when 16#0AA3# => romdata <= X"8610E028";
    when 16#0AA4# => romdata <= X"E400E008";
    when 16#0AA5# => romdata <= X"80A0C012";
    when 16#0AA6# => romdata <= X"2280002A";
    when 16#0AA7# => romdata <= X"C2046004";
    when 16#0AA8# => romdata <= X"C404A004";
    when 16#0AA9# => romdata <= X"8408BFFC";
    when 16#0AAA# => romdata <= X"82208010";
    when 16#0AAB# => romdata <= X"80A0600F";
    when 16#0AAC# => romdata <= X"1480008A";
    when 16#0AAD# => romdata <= X"80A06000";
    when 16#0AAE# => romdata <= X"C620E00C";
    when 16#0AAF# => romdata <= X"16800059";
    when 16#0AB0# => romdata <= X"C620E008";
    when 16#0AB1# => romdata <= X"80A0A1FF";
    when 16#0AB2# => romdata <= X"28800062";
    when 16#0AB3# => romdata <= X"8530A003";
    when 16#0AB4# => romdata <= X"8330A009";
    when 16#0AB5# => romdata <= X"80A06004";
    when 16#0AB6# => romdata <= X"188000E9";
    when 16#0AB7# => romdata <= X"8800605B";
    when 16#0AB8# => romdata <= X"8930A006";
    when 16#0AB9# => romdata <= X"88012038";
    when 16#0ABA# => romdata <= X"9B292003";
    when 16#0ABB# => romdata <= X"9A04400D";
    when 16#0ABC# => romdata <= X"C2036008";
    when 16#0ABD# => romdata <= X"80A0400D";
    when 16#0ABE# => romdata <= X"32800008";
    when 16#0ABF# => romdata <= X"C8006004";
    when 16#0AC0# => romdata <= X"108000E9";
    when 16#0AC1# => romdata <= X"DA046004";
    when 16#0AC2# => romdata <= X"80A34001";
    when 16#0AC3# => romdata <= X"22800008";
    when 16#0AC4# => romdata <= X"C400600C";
    when 16#0AC5# => romdata <= X"C8006004";
    when 16#0AC6# => romdata <= X"88093FFC";
    when 16#0AC7# => romdata <= X"80A08004";
    when 16#0AC8# => romdata <= X"2ABFFFFA";
    when 16#0AC9# => romdata <= X"C2006008";
    when 16#0ACA# => romdata <= X"C400600C";
    when 16#0ACB# => romdata <= X"C424A00C";
    when 16#0ACC# => romdata <= X"C224A008";
    when 16#0ACD# => romdata <= X"E420600C";
    when 16#0ACE# => romdata <= X"E420A008";
    when 16#0ACF# => romdata <= X"C2046004";
    when 16#0AD0# => romdata <= X"853B2002";
    when 16#0AD1# => romdata <= X"88102001";
    when 16#0AD2# => romdata <= X"89290002";
    when 16#0AD3# => romdata <= X"80A04004";
    when 16#0AD4# => romdata <= X"2ABFFF7E";
    when 16#0AD5# => romdata <= X"E6046008";
    when 16#0AD6# => romdata <= X"80884004";
    when 16#0AD7# => romdata <= X"2280004B";
    when 16#0AD8# => romdata <= X"980B3FFC";
    when 16#0AD9# => romdata <= X"952B2003";
    when 16#0ADA# => romdata <= X"9610000C";
    when 16#0ADB# => romdata <= X"9404400A";
    when 16#0ADC# => romdata <= X"9A10000A";
    when 16#0ADD# => romdata <= X"E403600C";
    when 16#0ADE# => romdata <= X"80A34012";
    when 16#0ADF# => romdata <= X"3280000B";
    when 16#0AE0# => romdata <= X"C404A004";
    when 16#0AE1# => romdata <= X"10800058";
    when 16#0AE2# => romdata <= X"9602E001";
    when 16#0AE3# => romdata <= X"36800019";
    when 16#0AE4# => romdata <= X"C604A00C";
    when 16#0AE5# => romdata <= X"E404A00C";
    when 16#0AE6# => romdata <= X"80A34012";
    when 16#0AE7# => romdata <= X"22800052";
    when 16#0AE8# => romdata <= X"9602E001";
    when 16#0AE9# => romdata <= X"C404A004";
    when 16#0AEA# => romdata <= X"8408BFFC";
    when 16#0AEB# => romdata <= X"82208010";
    when 16#0AEC# => romdata <= X"80A0600F";
    when 16#0AED# => romdata <= X"04BFFFF6";
    when 16#0AEE# => romdata <= X"80A06000";
    when 16#0AEF# => romdata <= X"DA04A00C";
    when 16#0AF0# => romdata <= X"C804A008";
    when 16#0AF1# => romdata <= X"84048010";
    when 16#0AF2# => romdata <= X"A0142001";
    when 16#0AF3# => romdata <= X"C8236008";
    when 16#0AF4# => romdata <= X"DA21200C";
    when 16#0AF5# => romdata <= X"C420E00C";
    when 16#0AF6# => romdata <= X"C420E008";
    when 16#0AF7# => romdata <= X"E024A004";
    when 16#0AF8# => romdata <= X"C2208001";
    when 16#0AF9# => romdata <= X"C620A008";
    when 16#0AFA# => romdata <= X"10800010";
    when 16#0AFB# => romdata <= X"C620A00C";
    when 16#0AFC# => romdata <= X"C204A008";
    when 16#0AFD# => romdata <= X"84048002";
    when 16#0AFE# => romdata <= X"C800A004";
    when 16#0AFF# => romdata <= X"88112001";
    when 16#0B00# => romdata <= X"C220E008";
    when 16#0B01# => romdata <= X"C820A004";
    when 16#0B02# => romdata <= X"C620600C";
    when 16#0B03# => romdata <= X"90100018";
    when 16#0B04# => romdata <= X"400000DB";
    when 16#0B05# => romdata <= X"B004A008";
    when 16#0B06# => romdata <= X"81C7E008";
    when 16#0B07# => romdata <= X"81E80000";
    when 16#0B08# => romdata <= X"84048002";
    when 16#0B09# => romdata <= X"C200A004";
    when 16#0B0A# => romdata <= X"82106001";
    when 16#0B0B# => romdata <= X"C220A004";
    when 16#0B0C# => romdata <= X"90100018";
    when 16#0B0D# => romdata <= X"400000D2";
    when 16#0B0E# => romdata <= X"B004A008";
    when 16#0B0F# => romdata <= X"81C7E008";
    when 16#0B10# => romdata <= X"81E80000";
    when 16#0B11# => romdata <= X"98032038";
    when 16#0B12# => romdata <= X"10BFFF79";
    when 16#0B13# => romdata <= X"872B2003";
    when 16#0B14# => romdata <= X"8928A003";
    when 16#0B15# => romdata <= X"88044004";
    when 16#0B16# => romdata <= X"DA012008";
    when 16#0B17# => romdata <= X"D6046004";
    when 16#0B18# => romdata <= X"C824A00C";
    when 16#0B19# => romdata <= X"DA24A008";
    when 16#0B1A# => romdata <= X"8538A002";
    when 16#0B1B# => romdata <= X"82102001";
    when 16#0B1C# => romdata <= X"E423600C";
    when 16#0B1D# => romdata <= X"83284002";
    when 16#0B1E# => romdata <= X"E4212008";
    when 16#0B1F# => romdata <= X"8210400B";
    when 16#0B20# => romdata <= X"10BFFFB0";
    when 16#0B21# => romdata <= X"C2246004";
    when 16#0B22# => romdata <= X"89292001";
    when 16#0B23# => romdata <= X"80884004";
    when 16#0B24# => romdata <= X"02BFFFFE";
    when 16#0B25# => romdata <= X"98032004";
    when 16#0B26# => romdata <= X"10BFFFB4";
    when 16#0B27# => romdata <= X"952B2003";
    when 16#0B28# => romdata <= X"38BFFF31";
    when 16#0B29# => romdata <= X"03100037";
    when 16#0B2A# => romdata <= X"E4046008";
    when 16#0B2B# => romdata <= X"84048010";
    when 16#0B2C# => romdata <= X"A0142001";
    when 16#0B2D# => romdata <= X"82106001";
    when 16#0B2E# => romdata <= X"E024A004";
    when 16#0B2F# => romdata <= X"C220A004";
    when 16#0B30# => romdata <= X"90100018";
    when 16#0B31# => romdata <= X"C4246008";
    when 16#0B32# => romdata <= X"400000AD";
    when 16#0B33# => romdata <= X"B004A008";
    when 16#0B34# => romdata <= X"81C7E008";
    when 16#0B35# => romdata <= X"81E80000";
    when 16#0B36# => romdata <= X"84048010";
    when 16#0B37# => romdata <= X"10BFFFBE";
    when 16#0B38# => romdata <= X"A0142001";
    when 16#0B39# => romdata <= X"808AE003";
    when 16#0B3A# => romdata <= X"12BFFFA3";
    when 16#0B3B# => romdata <= X"9A04A008";
    when 16#0B3C# => romdata <= X"808B2003";
    when 16#0B3D# => romdata <= X"0280009C";
    when 16#0B3E# => romdata <= X"8202BFF8";
    when 16#0B3F# => romdata <= X"D4006008";
    when 16#0B40# => romdata <= X"80A28001";
    when 16#0B41# => romdata <= X"22BFFFFB";
    when 16#0B42# => romdata <= X"98033FFF";
    when 16#0B43# => romdata <= X"C2046004";
    when 16#0B44# => romdata <= X"89292001";
    when 16#0B45# => romdata <= X"80A10001";
    when 16#0B46# => romdata <= X"18BFFF0B";
    when 16#0B47# => romdata <= X"80A12000";
    when 16#0B48# => romdata <= X"22BFFF0A";
    when 16#0B49# => romdata <= X"E6046008";
    when 16#0B4A# => romdata <= X"80890001";
    when 16#0B4B# => romdata <= X"22800092";
    when 16#0B4C# => romdata <= X"89292001";
    when 16#0B4D# => romdata <= X"10BFFF8C";
    when 16#0B4E# => romdata <= X"9810000B";
    when 16#0B4F# => romdata <= X"8204A008";
    when 16#0B50# => romdata <= X"E400600C";
    when 16#0B51# => romdata <= X"80A04012";
    when 16#0B52# => romdata <= X"02BFFF50";
    when 16#0B53# => romdata <= X"98032002";
    when 16#0B54# => romdata <= X"10BFFEEF";
    when 16#0B55# => romdata <= X"C604A004";
    when 16#0B56# => romdata <= X"C205A2FC";
    when 16#0B57# => romdata <= X"82054001";
    when 16#0B58# => romdata <= X"80A08012";
    when 16#0B59# => romdata <= X"02800067";
    when 16#0B5A# => romdata <= X"C225A2FC";
    when 16#0B5B# => romdata <= X"C605E02C";
    when 16#0B5C# => romdata <= X"80A0FFFF";
    when 16#0B5D# => romdata <= X"2280006B";
    when 16#0B5E# => romdata <= X"03100035";
    when 16#0B5F# => romdata <= X"82048001";
    when 16#0B60# => romdata <= X"84204002";
    when 16#0B61# => romdata <= X"C425A2FC";
    when 16#0B62# => romdata <= X"848CA007";
    when 16#0B63# => romdata <= X"02800006";
    when 16#0B64# => romdata <= X"03000004";
    when 16#0B65# => romdata <= X"82102008";
    when 16#0B66# => romdata <= X"82204002";
    when 16#0B67# => romdata <= X"A4048001";
    when 16#0B68# => romdata <= X"82207000";
    when 16#0B69# => romdata <= X"AA048015";
    when 16#0B6A# => romdata <= X"90100018";
    when 16#0B6B# => romdata <= X"AA0D6FFF";
    when 16#0B6C# => romdata <= X"AA204015";
    when 16#0B6D# => romdata <= X"4000007E";
    when 16#0B6E# => romdata <= X"92100015";
    when 16#0B6F# => romdata <= X"80A23FFF";
    when 16#0B70# => romdata <= X"02800060";
    when 16#0B71# => romdata <= X"84102001";
    when 16#0B72# => romdata <= X"84220012";
    when 16#0B73# => romdata <= X"84008015";
    when 16#0B74# => romdata <= X"8410A001";
    when 16#0B75# => romdata <= X"C205A2FC";
    when 16#0B76# => romdata <= X"82054001";
    when 16#0B77# => romdata <= X"C225A2FC";
    when 16#0B78# => romdata <= X"C424A004";
    when 16#0B79# => romdata <= X"80A44013";
    when 16#0B7A# => romdata <= X"02800010";
    when 16#0B7B# => romdata <= X"E4246008";
    when 16#0B7C# => romdata <= X"80A5200F";
    when 16#0B7D# => romdata <= X"0880003A";
    when 16#0B7E# => romdata <= X"84053FF4";
    when 16#0B7F# => romdata <= X"8408BFF8";
    when 16#0B80# => romdata <= X"8604C002";
    when 16#0B81# => romdata <= X"C804E004";
    when 16#0B82# => romdata <= X"88092001";
    when 16#0B83# => romdata <= X"88108004";
    when 16#0B84# => romdata <= X"C824E004";
    when 16#0B85# => romdata <= X"88102005";
    when 16#0B86# => romdata <= X"C820E008";
    when 16#0B87# => romdata <= X"80A0A00F";
    when 16#0B88# => romdata <= X"18800042";
    when 16#0B89# => romdata <= X"C820E004";
    when 16#0B8A# => romdata <= X"05100037";
    when 16#0B8B# => romdata <= X"C600A2F4";
    when 16#0B8C# => romdata <= X"80A04003";
    when 16#0B8D# => romdata <= X"38800002";
    when 16#0B8E# => romdata <= X"C220A2F4";
    when 16#0B8F# => romdata <= X"05100037";
    when 16#0B90# => romdata <= X"C600A2F8";
    when 16#0B91# => romdata <= X"80A04003";
    when 16#0B92# => romdata <= X"38BFFEDD";
    when 16#0B93# => romdata <= X"C220A2F8";
    when 16#0B94# => romdata <= X"10BFFEDC";
    when 16#0B95# => romdata <= X"C2046008";
    when 16#0B96# => romdata <= X"28BFFF95";
    when 16#0B97# => romdata <= X"E4046008";
    when 16#0B98# => romdata <= X"30BFFEDE";
    when 16#0B99# => romdata <= X"18800017";
    when 16#0B9A# => romdata <= X"80A06554";
    when 16#0B9B# => romdata <= X"9934200F";
    when 16#0B9C# => romdata <= X"98032077";
    when 16#0B9D# => romdata <= X"10BFFEEE";
    when 16#0B9E# => romdata <= X"872B2003";
    when 16#0B9F# => romdata <= X"80A06014";
    when 16#0BA0# => romdata <= X"08BFFF1B";
    when 16#0BA1# => romdata <= X"9B292003";
    when 16#0BA2# => romdata <= X"80A06054";
    when 16#0BA3# => romdata <= X"18800017";
    when 16#0BA4# => romdata <= X"80A06154";
    when 16#0BA5# => romdata <= X"8930A00C";
    when 16#0BA6# => romdata <= X"8801206E";
    when 16#0BA7# => romdata <= X"10BFFF14";
    when 16#0BA8# => romdata <= X"9B292003";
    when 16#0BA9# => romdata <= X"89392002";
    when 16#0BAA# => romdata <= X"84102001";
    when 16#0BAB# => romdata <= X"85288004";
    when 16#0BAC# => romdata <= X"84134002";
    when 16#0BAD# => romdata <= X"C4246004";
    when 16#0BAE# => romdata <= X"10BFFF1D";
    when 16#0BAF# => romdata <= X"84100001";
    when 16#0BB0# => romdata <= X"861023F0";
    when 16#0BB1# => romdata <= X"18BFFEDA";
    when 16#0BB2# => romdata <= X"9810207E";
    when 16#0BB3# => romdata <= X"99342012";
    when 16#0BB4# => romdata <= X"9803207C";
    when 16#0BB5# => romdata <= X"10BFFED6";
    when 16#0BB6# => romdata <= X"872B2003";
    when 16#0BB7# => romdata <= X"82102001";
    when 16#0BB8# => romdata <= X"10BFFEB7";
    when 16#0BB9# => romdata <= X"C224A004";
    when 16#0BBA# => romdata <= X"18800018";
    when 16#0BBB# => romdata <= X"80A06554";
    when 16#0BBC# => romdata <= X"8930A00F";
    when 16#0BBD# => romdata <= X"88012077";
    when 16#0BBE# => romdata <= X"10BFFEFD";
    when 16#0BBF# => romdata <= X"9B292003";
    when 16#0BC0# => romdata <= X"8088AFFF";
    when 16#0BC1# => romdata <= X"12BFFF9B";
    when 16#0BC2# => romdata <= X"C605E02C";
    when 16#0BC3# => romdata <= X"C4046008";
    when 16#0BC4# => romdata <= X"86054014";
    when 16#0BC5# => romdata <= X"8610E001";
    when 16#0BC6# => romdata <= X"10BFFFC4";
    when 16#0BC7# => romdata <= X"C620A004";
    when 16#0BC8# => romdata <= X"10BFFF9A";
    when 16#0BC9# => romdata <= X"E420602C";
    when 16#0BCA# => romdata <= X"9204E008";
    when 16#0BCB# => romdata <= X"4000106C";
    when 16#0BCC# => romdata <= X"90100018";
    when 16#0BCD# => romdata <= X"03100037";
    when 16#0BCE# => romdata <= X"10BFFFBC";
    when 16#0BCF# => romdata <= X"C20062FC";
    when 16#0BD0# => romdata <= X"10BFFFA5";
    when 16#0BD1# => romdata <= X"AA102000";
    when 16#0BD2# => romdata <= X"9A1023F0";
    when 16#0BD3# => romdata <= X"18BFFEE8";
    when 16#0BD4# => romdata <= X"8810207E";
    when 16#0BD5# => romdata <= X"8930A012";
    when 16#0BD6# => romdata <= X"8801207C";
    when 16#0BD7# => romdata <= X"10BFFEE4";
    when 16#0BD8# => romdata <= X"9B292003";
    when 16#0BD9# => romdata <= X"C2046004";
    when 16#0BDA# => romdata <= X"82284004";
    when 16#0BDB# => romdata <= X"10BFFF68";
    when 16#0BDC# => romdata <= X"C2246004";
    when 16#0BDD# => romdata <= X"10BFFF6D";
    when 16#0BDE# => romdata <= X"9602E004";
    when 16#0BDF# => romdata <= X"11100035";
    when 16#0BE0# => romdata <= X"90122030";
    when 16#0BE1# => romdata <= X"8213C000";
    when 16#0BE2# => romdata <= X"40001ED8";
    when 16#0BE3# => romdata <= X"9E104000";
    when 16#0BE4# => romdata <= X"01000000";
    when 16#0BE5# => romdata <= X"11100035";
    when 16#0BE6# => romdata <= X"90122030";
    when 16#0BE7# => romdata <= X"8213C000";
    when 16#0BE8# => romdata <= X"40001EBC";
    when 16#0BE9# => romdata <= X"9E104000";
    when 16#0BEA# => romdata <= X"01000000";
    when 16#0BEB# => romdata <= X"9DE3BFA0";
    when 16#0BEC# => romdata <= X"21100038";
    when 16#0BED# => romdata <= X"90100019";
    when 16#0BEE# => romdata <= X"40001C59";
    when 16#0BEF# => romdata <= X"C0242260";
    when 16#0BF0# => romdata <= X"80A23FFF";
    when 16#0BF1# => romdata <= X"02800004";
    when 16#0BF2# => romdata <= X"C2042260";
    when 16#0BF3# => romdata <= X"81C7E008";
    when 16#0BF4# => romdata <= X"91E80008";
    when 16#0BF5# => romdata <= X"80A06000";
    when 16#0BF6# => romdata <= X"02BFFFFD";
    when 16#0BF7# => romdata <= X"01000000";
    when 16#0BF8# => romdata <= X"C2260000";
    when 16#0BF9# => romdata <= X"81C7E008";
    when 16#0BFA# => romdata <= X"91E80008";
    when 16#0BFB# => romdata <= X"40004228";
    when 16#0BFC# => romdata <= X"400032FC";
    when 16#0BFD# => romdata <= X"400032FC";
    when 16#0BFE# => romdata <= X"4000400C";
    when 16#0BFF# => romdata <= X"400032FC";
    when 16#0C00# => romdata <= X"400032FC";
    when 16#0C01# => romdata <= X"400032FC";
    when 16#0C02# => romdata <= X"400032FC";
    when 16#0C03# => romdata <= X"400032FC";
    when 16#0C04# => romdata <= X"400032FC";
    when 16#0C05# => romdata <= X"40003F7C";
    when 16#0C06# => romdata <= X"40004028";
    when 16#0C07# => romdata <= X"400032FC";
    when 16#0C08# => romdata <= X"40003F90";
    when 16#0C09# => romdata <= X"4000412C";
    when 16#0C0A# => romdata <= X"400032FC";
    when 16#0C0B# => romdata <= X"40004038";
    when 16#0C0C# => romdata <= X"40004048";
    when 16#0C0D# => romdata <= X"40004048";
    when 16#0C0E# => romdata <= X"40004048";
    when 16#0C0F# => romdata <= X"40004048";
    when 16#0C10# => romdata <= X"40004048";
    when 16#0C11# => romdata <= X"40004048";
    when 16#0C12# => romdata <= X"40004048";
    when 16#0C13# => romdata <= X"40004048";
    when 16#0C14# => romdata <= X"40004048";
    when 16#0C15# => romdata <= X"400032FC";
    when 16#0C16# => romdata <= X"400032FC";
    when 16#0C17# => romdata <= X"400032FC";
    when 16#0C18# => romdata <= X"400032FC";
    when 16#0C19# => romdata <= X"400032FC";
    when 16#0C1A# => romdata <= X"400032FC";
    when 16#0C1B# => romdata <= X"400032FC";
    when 16#0C1C# => romdata <= X"400032FC";
    when 16#0C1D# => romdata <= X"400032FC";
    when 16#0C1E# => romdata <= X"40003FA0";
    when 16#0C1F# => romdata <= X"4000370C";
    when 16#0C20# => romdata <= X"40004258";
    when 16#0C21# => romdata <= X"400032FC";
    when 16#0C22# => romdata <= X"40004258";
    when 16#0C23# => romdata <= X"400032FC";
    when 16#0C24# => romdata <= X"400032FC";
    when 16#0C25# => romdata <= X"400032FC";
    when 16#0C26# => romdata <= X"400032FC";
    when 16#0C27# => romdata <= X"40004248";
    when 16#0C28# => romdata <= X"400032FC";
    when 16#0C29# => romdata <= X"400032FC";
    when 16#0C2A# => romdata <= X"400036C4";
    when 16#0C2B# => romdata <= X"400032FC";
    when 16#0C2C# => romdata <= X"400032FC";
    when 16#0C2D# => romdata <= X"400032FC";
    when 16#0C2E# => romdata <= X"40004198";
    when 16#0C2F# => romdata <= X"400032FC";
    when 16#0C30# => romdata <= X"400035F4";
    when 16#0C31# => romdata <= X"400032FC";
    when 16#0C32# => romdata <= X"400032FC";
    when 16#0C33# => romdata <= X"40004208";
    when 16#0C34# => romdata <= X"400032FC";
    when 16#0C35# => romdata <= X"400032FC";
    when 16#0C36# => romdata <= X"400032FC";
    when 16#0C37# => romdata <= X"400032FC";
    when 16#0C38# => romdata <= X"400032FC";
    when 16#0C39# => romdata <= X"400032FC";
    when 16#0C3A# => romdata <= X"400032FC";
    when 16#0C3B# => romdata <= X"400032FC";
    when 16#0C3C# => romdata <= X"400032FC";
    when 16#0C3D# => romdata <= X"400032FC";
    when 16#0C3E# => romdata <= X"40003FA0";
    when 16#0C3F# => romdata <= X"40003710";
    when 16#0C40# => romdata <= X"40004258";
    when 16#0C41# => romdata <= X"40004258";
    when 16#0C42# => romdata <= X"40004258";
    when 16#0C43# => romdata <= X"40004188";
    when 16#0C44# => romdata <= X"40003710";
    when 16#0C45# => romdata <= X"400032FC";
    when 16#0C46# => romdata <= X"400032FC";
    when 16#0C47# => romdata <= X"400040B8";
    when 16#0C48# => romdata <= X"400032FC";
    when 16#0C49# => romdata <= X"40003FE8";
    when 16#0C4A# => romdata <= X"400036C8";
    when 16#0C4B# => romdata <= X"4000407C";
    when 16#0C4C# => romdata <= X"400040A8";
    when 16#0C4D# => romdata <= X"400032FC";
    when 16#0C4E# => romdata <= X"40004198";
    when 16#0C4F# => romdata <= X"400032FC";
    when 16#0C50# => romdata <= X"400035F8";
    when 16#0C51# => romdata <= X"400032FC";
    when 16#0C52# => romdata <= X"400032FC";
    when 16#0C53# => romdata <= X"400040D8";
    when 16#0C54# => romdata <= X"9DE3BFA0";
    when 16#0C55# => romdata <= X"C2066008";
    when 16#0C56# => romdata <= X"80A06000";
    when 16#0C57# => romdata <= X"12800005";
    when 16#0C58# => romdata <= X"90100018";
    when 16#0C59# => romdata <= X"C0266004";
    when 16#0C5A# => romdata <= X"81C7E008";
    when 16#0C5B# => romdata <= X"91E82000";
    when 16#0C5C# => romdata <= X"40001082";
    when 16#0C5D# => romdata <= X"92100019";
    when 16#0C5E# => romdata <= X"C0266004";
    when 16#0C5F# => romdata <= X"C0266008";
    when 16#0C60# => romdata <= X"81C7E008";
    when 16#0C61# => romdata <= X"91E80008";
    when 16#0C62# => romdata <= X"9DE3B870";
    when 16#0C63# => romdata <= X"400011FA";
    when 16#0C64# => romdata <= X"01000000";
    when 16#0C65# => romdata <= X"D0020000";
    when 16#0C66# => romdata <= X"C216600C";
    when 16#0C67# => romdata <= X"F027A044";
    when 16#0C68# => romdata <= X"80886200";
    when 16#0C69# => romdata <= X"02800308";
    when 16#0C6A# => romdata <= X"D027B8E8";
    when 16#0C6B# => romdata <= X"03100032";
    when 16#0C6C# => romdata <= X"D00062C8";
    when 16#0C6D# => romdata <= X"80A22000";
    when 16#0C6E# => romdata <= X"22800007";
    when 16#0C6F# => romdata <= X"C216600C";
    when 16#0C70# => romdata <= X"C2022038";
    when 16#0C71# => romdata <= X"80A06000";
    when 16#0C72# => romdata <= X"02800303";
    when 16#0C73# => romdata <= X"01000000";
    when 16#0C74# => romdata <= X"C216600C";
    when 16#0C75# => romdata <= X"80886008";
    when 16#0C76# => romdata <= X"0280026E";
    when 16#0C77# => romdata <= X"86100001";
    when 16#0C78# => romdata <= X"C4066010";
    when 16#0C79# => romdata <= X"80A0A000";
    when 16#0C7A# => romdata <= X"0280026A";
    when 16#0C7B# => romdata <= X"8408601A";
    when 16#0C7C# => romdata <= X"80A0A00A";
    when 16#0C7D# => romdata <= X"22800273";
    when 16#0C7E# => romdata <= X"C456600E";
    when 16#0C7F# => romdata <= X"A607BF40";
    when 16#0C80# => romdata <= X"C027BFB4";
    when 16#0C81# => romdata <= X"C027BFB0";
    when 16#0C82# => romdata <= X"E627BFAC";
    when 16#0C83# => romdata <= X"C027B8F8";
    when 16#0C84# => romdata <= X"C027B8FC";
    when 16#0C85# => romdata <= X"C027B8EC";
    when 16#0C86# => romdata <= X"C027B8F0";
    when 16#0C87# => romdata <= X"25100032";
    when 16#0C88# => romdata <= X"23100032";
    when 16#0C89# => romdata <= X"A414A078";
    when 16#0C8A# => romdata <= X"A2146068";
    when 16#0C8B# => romdata <= X"B0102000";
    when 16#0C8C# => romdata <= X"A0100013";
    when 16#0C8D# => romdata <= X"C44E8000";
    when 16#0C8E# => romdata <= X"80A0A025";
    when 16#0C8F# => romdata <= X"0280001E";
    when 16#0C90# => romdata <= X"C20E8000";
    when 16#0C91# => romdata <= X"80A0A000";
    when 16#0C92# => romdata <= X"0280001C";
    when 16#0C93# => romdata <= X"83286018";
    when 16#0C94# => romdata <= X"A810001A";
    when 16#0C95# => romdata <= X"A8052001";
    when 16#0C96# => romdata <= X"C24D0000";
    when 16#0C97# => romdata <= X"80A06025";
    when 16#0C98# => romdata <= X"02800004";
    when 16#0C99# => romdata <= X"80A06000";
    when 16#0C9A# => romdata <= X"32BFFFFC";
    when 16#0C9B# => romdata <= X"A8052001";
    when 16#0C9C# => romdata <= X"AAA5001A";
    when 16#0C9D# => romdata <= X"228000DE";
    when 16#0C9E# => romdata <= X"B4100014";
    when 16#0C9F# => romdata <= X"EA242004";
    when 16#0CA0# => romdata <= X"F4240000";
    when 16#0CA1# => romdata <= X"A0042008";
    when 16#0CA2# => romdata <= X"C207BFB0";
    when 16#0CA3# => romdata <= X"C407BFB4";
    when 16#0CA4# => romdata <= X"82006001";
    when 16#0CA5# => romdata <= X"84008015";
    when 16#0CA6# => romdata <= X"C227BFB0";
    when 16#0CA7# => romdata <= X"80A06007";
    when 16#0CA8# => romdata <= X"148002C1";
    when 16#0CA9# => romdata <= X"C427BFB4";
    when 16#0CAA# => romdata <= X"C20D0000";
    when 16#0CAB# => romdata <= X"B4100014";
    when 16#0CAC# => romdata <= X"B0060015";
    when 16#0CAD# => romdata <= X"83286018";
    when 16#0CAE# => romdata <= X"80A06000";
    when 16#0CAF# => romdata <= X"02800576";
    when 16#0CB0# => romdata <= X"B406A001";
    when 16#0CB1# => romdata <= X"C02FBFFF";
    when 16#0CB2# => romdata <= X"AC103FFF";
    when 16#0CB3# => romdata <= X"EA0E8000";
    when 16#0CB4# => romdata <= X"AB2D6018";
    when 16#0CB5# => romdata <= X"B8102000";
    when 16#0CB6# => romdata <= X"A8102000";
    when 16#0CB7# => romdata <= X"8610202B";
    when 16#0CB8# => romdata <= X"88102020";
    when 16#0CB9# => romdata <= X"AB3D6018";
    when 16#0CBA# => romdata <= X"B406A001";
    when 16#0CBB# => romdata <= X"82057FE0";
    when 16#0CBC# => romdata <= X"80A06058";
    when 16#0CBD# => romdata <= X"288000B9";
    when 16#0CBE# => romdata <= X"83286002";
    when 16#0CBF# => romdata <= X"80A56000";
    when 16#0CC0# => romdata <= X"02800565";
    when 16#0CC1# => romdata <= X"84102001";
    when 16#0CC2# => romdata <= X"EA2FBD18";
    when 16#0CC3# => romdata <= X"C02FBFFF";
    when 16#0CC4# => romdata <= X"C427B910";
    when 16#0CC5# => romdata <= X"C027B908";
    when 16#0CC6# => romdata <= X"BA102001";
    when 16#0CC7# => romdata <= X"AE07BD18";
    when 16#0CC8# => romdata <= X"AC102000";
    when 16#0CC9# => romdata <= X"808D2002";
    when 16#0CCA# => romdata <= X"0280011A";
    when 16#0CCB# => romdata <= X"868D2084";
    when 16#0CCC# => romdata <= X"C407B910";
    when 16#0CCD# => romdata <= X"8400A002";
    when 16#0CCE# => romdata <= X"C427B910";
    when 16#0CCF# => romdata <= X"02800117";
    when 16#0CD0# => romdata <= X"C627B90C";
    when 16#0CD1# => romdata <= X"C24FBFFF";
    when 16#0CD2# => romdata <= X"80A06000";
    when 16#0CD3# => romdata <= X"02800152";
    when 16#0CD4# => romdata <= X"808D2002";
    when 16#0CD5# => romdata <= X"82102001";
    when 16#0CD6# => romdata <= X"C2242004";
    when 16#0CD7# => romdata <= X"8207BFFF";
    when 16#0CD8# => romdata <= X"C2240000";
    when 16#0CD9# => romdata <= X"C407BFB4";
    when 16#0CDA# => romdata <= X"C207BFB0";
    when 16#0CDB# => romdata <= X"82006001";
    when 16#0CDC# => romdata <= X"8400A001";
    when 16#0CDD# => romdata <= X"C227BFB0";
    when 16#0CDE# => romdata <= X"C427BFB4";
    when 16#0CDF# => romdata <= X"80A06007";
    when 16#0CE0# => romdata <= X"14800157";
    when 16#0CE1# => romdata <= X"A0042008";
    when 16#0CE2# => romdata <= X"C207B90C";
    when 16#0CE3# => romdata <= X"80A06080";
    when 16#0CE4# => romdata <= X"0280015D";
    when 16#0CE5# => romdata <= X"C407B910";
    when 16#0CE6# => romdata <= X"C407B908";
    when 16#0CE7# => romdata <= X"8220801D";
    when 16#0CE8# => romdata <= X"80A06000";
    when 16#0CE9# => romdata <= X"04800038";
    when 16#0CEA# => romdata <= X"80A06010";
    when 16#0CEB# => romdata <= X"04800024";
    when 16#0CEC# => romdata <= X"E227B90C";
    when 16#0CED# => romdata <= X"86100010";
    when 16#0CEE# => romdata <= X"84102010";
    when 16#0CEF# => romdata <= X"A0100001";
    when 16#0CF0# => romdata <= X"10800006";
    when 16#0CF1# => romdata <= X"82100003";
    when 16#0CF2# => romdata <= X"A0043FF0";
    when 16#0CF3# => romdata <= X"80A42010";
    when 16#0CF4# => romdata <= X"24800019";
    when 16#0CF5# => romdata <= X"84100001";
    when 16#0CF6# => romdata <= X"C4206004";
    when 16#0CF7# => romdata <= X"E2204000";
    when 16#0CF8# => romdata <= X"82006008";
    when 16#0CF9# => romdata <= X"C607BFB0";
    when 16#0CFA# => romdata <= X"C807BFB4";
    when 16#0CFB# => romdata <= X"8600E001";
    when 16#0CFC# => romdata <= X"88012010";
    when 16#0CFD# => romdata <= X"C627BFB0";
    when 16#0CFE# => romdata <= X"80A0E007";
    when 16#0CFF# => romdata <= X"04BFFFF3";
    when 16#0D00# => romdata <= X"C827BFB4";
    when 16#0D01# => romdata <= X"C427B8E4";
    when 16#0D02# => romdata <= X"90100019";
    when 16#0D03# => romdata <= X"7FFFFF51";
    when 16#0D04# => romdata <= X"9207BFAC";
    when 16#0D05# => romdata <= X"80A22000";
    when 16#0D06# => romdata <= X"128001CB";
    when 16#0D07# => romdata <= X"C407B8E4";
    when 16#0D08# => romdata <= X"A0043FF0";
    when 16#0D09# => romdata <= X"80A42010";
    when 16#0D0A# => romdata <= X"14BFFFEC";
    when 16#0D0B# => romdata <= X"82100013";
    when 16#0D0C# => romdata <= X"84100001";
    when 16#0D0D# => romdata <= X"82100010";
    when 16#0D0E# => romdata <= X"A0100002";
    when 16#0D0F# => romdata <= X"C2242004";
    when 16#0D10# => romdata <= X"C607B90C";
    when 16#0D11# => romdata <= X"C6240000";
    when 16#0D12# => romdata <= X"C407BFB4";
    when 16#0D13# => romdata <= X"82008001";
    when 16#0D14# => romdata <= X"C227BFB4";
    when 16#0D15# => romdata <= X"C207BFB0";
    when 16#0D16# => romdata <= X"82006001";
    when 16#0D17# => romdata <= X"C227BFB0";
    when 16#0D18# => romdata <= X"80A06007";
    when 16#0D19# => romdata <= X"04800008";
    when 16#0D1A# => romdata <= X"A0042008";
    when 16#0D1B# => romdata <= X"90100019";
    when 16#0D1C# => romdata <= X"7FFFFF38";
    when 16#0D1D# => romdata <= X"9207BFAC";
    when 16#0D1E# => romdata <= X"80A22000";
    when 16#0D1F# => romdata <= X"128001B2";
    when 16#0D20# => romdata <= X"A0100013";
    when 16#0D21# => romdata <= X"808D2100";
    when 16#0D22# => romdata <= X"1280015B";
    when 16#0D23# => romdata <= X"80A56065";
    when 16#0D24# => romdata <= X"FA242004";
    when 16#0D25# => romdata <= X"EE240000";
    when 16#0D26# => romdata <= X"A0042008";
    when 16#0D27# => romdata <= X"C207BFB4";
    when 16#0D28# => romdata <= X"BA00401D";
    when 16#0D29# => romdata <= X"FA27BFB4";
    when 16#0D2A# => romdata <= X"C207BFB0";
    when 16#0D2B# => romdata <= X"82006001";
    when 16#0D2C# => romdata <= X"80A06007";
    when 16#0D2D# => romdata <= X"14800234";
    when 16#0D2E# => romdata <= X"C227BFB0";
    when 16#0D2F# => romdata <= X"808D2004";
    when 16#0D30# => romdata <= X"02800036";
    when 16#0D31# => romdata <= X"E807BFB4";
    when 16#0D32# => romdata <= X"C207B910";
    when 16#0D33# => romdata <= X"A8270001";
    when 16#0D34# => romdata <= X"80A52000";
    when 16#0D35# => romdata <= X"04800030";
    when 16#0D36# => romdata <= X"80A52010";
    when 16#0D37# => romdata <= X"0480001D";
    when 16#0D38# => romdata <= X"E427B904";
    when 16#0D39# => romdata <= X"AA102010";
    when 16#0D3A# => romdata <= X"10800006";
    when 16#0D3B# => romdata <= X"AE07BFAC";
    when 16#0D3C# => romdata <= X"A8053FF0";
    when 16#0D3D# => romdata <= X"80A52010";
    when 16#0D3E# => romdata <= X"24800017";
    when 16#0D3F# => romdata <= X"E8242004";
    when 16#0D40# => romdata <= X"EA242004";
    when 16#0D41# => romdata <= X"E4240000";
    when 16#0D42# => romdata <= X"A0042008";
    when 16#0D43# => romdata <= X"C207BFB0";
    when 16#0D44# => romdata <= X"C407BFB4";
    when 16#0D45# => romdata <= X"82006001";
    when 16#0D46# => romdata <= X"8400A010";
    when 16#0D47# => romdata <= X"C227BFB0";
    when 16#0D48# => romdata <= X"80A06007";
    when 16#0D49# => romdata <= X"04BFFFF3";
    when 16#0D4A# => romdata <= X"C427BFB4";
    when 16#0D4B# => romdata <= X"90100019";
    when 16#0D4C# => romdata <= X"7FFFFF08";
    when 16#0D4D# => romdata <= X"92100017";
    when 16#0D4E# => romdata <= X"80A22000";
    when 16#0D4F# => romdata <= X"12800182";
    when 16#0D50# => romdata <= X"A8053FF0";
    when 16#0D51# => romdata <= X"80A52010";
    when 16#0D52# => romdata <= X"14BFFFEE";
    when 16#0D53# => romdata <= X"A0100013";
    when 16#0D54# => romdata <= X"E8242004";
    when 16#0D55# => romdata <= X"C407B904";
    when 16#0D56# => romdata <= X"C4240000";
    when 16#0D57# => romdata <= X"C207BFB4";
    when 16#0D58# => romdata <= X"A8050001";
    when 16#0D59# => romdata <= X"C207BFB0";
    when 16#0D5A# => romdata <= X"82006001";
    when 16#0D5B# => romdata <= X"E827BFB4";
    when 16#0D5C# => romdata <= X"80A06007";
    when 16#0D5D# => romdata <= X"04800009";
    when 16#0D5E# => romdata <= X"C227BFB0";
    when 16#0D5F# => romdata <= X"90100019";
    when 16#0D60# => romdata <= X"7FFFFEF4";
    when 16#0D61# => romdata <= X"9207BFAC";
    when 16#0D62# => romdata <= X"80A22000";
    when 16#0D63# => romdata <= X"1280016F";
    when 16#0D64# => romdata <= X"80A5A000";
    when 16#0D65# => romdata <= X"E807BFB4";
    when 16#0D66# => romdata <= X"C607B910";
    when 16#0D67# => romdata <= X"80A70003";
    when 16#0D68# => romdata <= X"26800002";
    when 16#0D69# => romdata <= X"B8100003";
    when 16#0D6A# => romdata <= X"80A52000";
    when 16#0D6B# => romdata <= X"12800160";
    when 16#0D6C# => romdata <= X"B006001C";
    when 16#0D6D# => romdata <= X"C027BFB0";
    when 16#0D6E# => romdata <= X"80A5A000";
    when 16#0D6F# => romdata <= X"02BFFF1E";
    when 16#0D70# => romdata <= X"A0100013";
    when 16#0D71# => romdata <= X"D007A044";
    when 16#0D72# => romdata <= X"40000EC5";
    when 16#0D73# => romdata <= X"92100016";
    when 16#0D74# => romdata <= X"10BFFF1A";
    when 16#0D75# => romdata <= X"C44E8000";
    when 16#0D76# => romdata <= X"0510000B";
    when 16#0D77# => romdata <= X"8410A3EC";
    when 16#0D78# => romdata <= X"C2008001";
    when 16#0D79# => romdata <= X"81C04000";
    when 16#0D7A# => romdata <= X"01000000";
    when 16#0D7B# => romdata <= X"10BFFF32";
    when 16#0D7C# => romdata <= X"C20D0000";
    when 16#0D7D# => romdata <= X"A8152010";
    when 16#0D7E# => romdata <= X"808D2010";
    when 16#0D7F# => romdata <= X"3280002D";
    when 16#0D80# => romdata <= X"FA06C000";
    when 16#0D81# => romdata <= X"808D2040";
    when 16#0D82# => romdata <= X"2280002A";
    when 16#0D83# => romdata <= X"FA06C000";
    when 16#0D84# => romdata <= X"FA16E002";
    when 16#0D85# => romdata <= X"80A0001D";
    when 16#0D86# => romdata <= X"B606E004";
    when 16#0D87# => romdata <= X"84402000";
    when 16#0D88# => romdata <= X"82102001";
    when 16#0D89# => romdata <= X"C02FBFFF";
    when 16#0D8A# => romdata <= X"80A5A000";
    when 16#0D8B# => romdata <= X"36800002";
    when 16#0D8C# => romdata <= X"A80D3F7F";
    when 16#0D8D# => romdata <= X"8607BE74";
    when 16#0D8E# => romdata <= X"80A5A000";
    when 16#0D8F# => romdata <= X"12800005";
    when 16#0D90# => romdata <= X"C627B8DC";
    when 16#0D91# => romdata <= X"8088A0FF";
    when 16#0D92# => romdata <= X"0280003D";
    when 16#0D93# => romdata <= X"808860FF";
    when 16#0D94# => romdata <= X"820860FF";
    when 16#0D95# => romdata <= X"80A06001";
    when 16#0D96# => romdata <= X"02800333";
    when 16#0D97# => romdata <= X"80A06002";
    when 16#0D98# => romdata <= X"02800326";
    when 16#0D99# => romdata <= X"AE07BE74";
    when 16#0D9A# => romdata <= X"820F6007";
    when 16#0D9B# => romdata <= X"AE05FFFF";
    when 16#0D9C# => romdata <= X"82006030";
    when 16#0D9D# => romdata <= X"BB376003";
    when 16#0D9E# => romdata <= X"80A76000";
    when 16#0D9F# => romdata <= X"12BFFFFB";
    when 16#0DA0# => romdata <= X"C22DC000";
    when 16#0DA1# => romdata <= X"C407B8DC";
    when 16#0DA2# => romdata <= X"808D2001";
    when 16#0DA3# => romdata <= X"02800033";
    when 16#0DA4# => romdata <= X"BA208017";
    when 16#0DA5# => romdata <= X"80A06030";
    when 16#0DA6# => romdata <= X"02800030";
    when 16#0DA7# => romdata <= X"82102030";
    when 16#0DA8# => romdata <= X"AE05FFFF";
    when 16#0DA9# => romdata <= X"BA208017";
    when 16#0DAA# => romdata <= X"1080002C";
    when 16#0DAB# => romdata <= X"C22DC000";
    when 16#0DAC# => romdata <= X"80A0001D";
    when 16#0DAD# => romdata <= X"B606E004";
    when 16#0DAE# => romdata <= X"84402000";
    when 16#0DAF# => romdata <= X"10BFFFDA";
    when 16#0DB0# => romdata <= X"82102001";
    when 16#0DB1# => romdata <= X"A8152010";
    when 16#0DB2# => romdata <= X"808D2010";
    when 16#0DB3# => romdata <= X"3280000B";
    when 16#0DB4# => romdata <= X"FA06C000";
    when 16#0DB5# => romdata <= X"808D2040";
    when 16#0DB6# => romdata <= X"22800008";
    when 16#0DB7# => romdata <= X"FA06C000";
    when 16#0DB8# => romdata <= X"FA16E002";
    when 16#0DB9# => romdata <= X"80A0001D";
    when 16#0DBA# => romdata <= X"B606E004";
    when 16#0DBB# => romdata <= X"84402000";
    when 16#0DBC# => romdata <= X"10BFFFCD";
    when 16#0DBD# => romdata <= X"82102000";
    when 16#0DBE# => romdata <= X"80A0001D";
    when 16#0DBF# => romdata <= X"B606E004";
    when 16#0DC0# => romdata <= X"84402000";
    when 16#0DC1# => romdata <= X"10BFFFC8";
    when 16#0DC2# => romdata <= X"82102000";
    when 16#0DC3# => romdata <= X"A8152010";
    when 16#0DC4# => romdata <= X"808D2010";
    when 16#0DC5# => romdata <= X"02800210";
    when 16#0DC6# => romdata <= X"808D2040";
    when 16#0DC7# => romdata <= X"FA06C000";
    when 16#0DC8# => romdata <= X"B606E004";
    when 16#0DC9# => romdata <= X"80A76000";
    when 16#0DCA# => romdata <= X"06800352";
    when 16#0DCB# => romdata <= X"80A0001D";
    when 16#0DCC# => romdata <= X"82102001";
    when 16#0DCD# => romdata <= X"10BFFFBD";
    when 16#0DCE# => romdata <= X"84402000";
    when 16#0DCF# => romdata <= X"12800006";
    when 16#0DD0# => romdata <= X"AE07BE74";
    when 16#0DD1# => romdata <= X"808D2001";
    when 16#0DD2# => romdata <= X"128001DF";
    when 16#0DD3# => romdata <= X"82102030";
    when 16#0DD4# => romdata <= X"AE07BE74";
    when 16#0DD5# => romdata <= X"BA102000";
    when 16#0DD6# => romdata <= X"80A74016";
    when 16#0DD7# => romdata <= X"16800003";
    when 16#0DD8# => romdata <= X"FA27B910";
    when 16#0DD9# => romdata <= X"EC27B910";
    when 16#0DDA# => romdata <= X"EC27B908";
    when 16#0DDB# => romdata <= X"AC102000";
    when 16#0DDC# => romdata <= X"C24FBFFF";
    when 16#0DDD# => romdata <= X"80A06000";
    when 16#0DDE# => romdata <= X"02BFFEEC";
    when 16#0DDF# => romdata <= X"808D2002";
    when 16#0DE0# => romdata <= X"C207B910";
    when 16#0DE1# => romdata <= X"82006001";
    when 16#0DE2# => romdata <= X"C227B910";
    when 16#0DE3# => romdata <= X"868D2084";
    when 16#0DE4# => romdata <= X"12BFFEED";
    when 16#0DE5# => romdata <= X"C627B90C";
    when 16#0DE6# => romdata <= X"C407B910";
    when 16#0DE7# => romdata <= X"82270002";
    when 16#0DE8# => romdata <= X"80A06000";
    when 16#0DE9# => romdata <= X"04BFFEE8";
    when 16#0DEA# => romdata <= X"80A06010";
    when 16#0DEB# => romdata <= X"04800024";
    when 16#0DEC# => romdata <= X"E427B904";
    when 16#0DED# => romdata <= X"86100010";
    when 16#0DEE# => romdata <= X"84102010";
    when 16#0DEF# => romdata <= X"A0100001";
    when 16#0DF0# => romdata <= X"10800006";
    when 16#0DF1# => romdata <= X"82100003";
    when 16#0DF2# => romdata <= X"A0043FF0";
    when 16#0DF3# => romdata <= X"80A42010";
    when 16#0DF4# => romdata <= X"24800019";
    when 16#0DF5# => romdata <= X"84100001";
    when 16#0DF6# => romdata <= X"C4206004";
    when 16#0DF7# => romdata <= X"E4204000";
    when 16#0DF8# => romdata <= X"82006008";
    when 16#0DF9# => romdata <= X"C607BFB0";
    when 16#0DFA# => romdata <= X"C807BFB4";
    when 16#0DFB# => romdata <= X"8600E001";
    when 16#0DFC# => romdata <= X"88012010";
    when 16#0DFD# => romdata <= X"C627BFB0";
    when 16#0DFE# => romdata <= X"80A0E007";
    when 16#0DFF# => romdata <= X"04BFFFF3";
    when 16#0E00# => romdata <= X"C827BFB4";
    when 16#0E01# => romdata <= X"C427B8E4";
    when 16#0E02# => romdata <= X"90100019";
    when 16#0E03# => romdata <= X"7FFFFE51";
    when 16#0E04# => romdata <= X"9207BFAC";
    when 16#0E05# => romdata <= X"80A22000";
    when 16#0E06# => romdata <= X"128000CB";
    when 16#0E07# => romdata <= X"C407B8E4";
    when 16#0E08# => romdata <= X"A0043FF0";
    when 16#0E09# => romdata <= X"80A42010";
    when 16#0E0A# => romdata <= X"14BFFFEC";
    when 16#0E0B# => romdata <= X"82100013";
    when 16#0E0C# => romdata <= X"84100001";
    when 16#0E0D# => romdata <= X"82100010";
    when 16#0E0E# => romdata <= X"A0100002";
    when 16#0E0F# => romdata <= X"C2242004";
    when 16#0E10# => romdata <= X"C607B904";
    when 16#0E11# => romdata <= X"C6240000";
    when 16#0E12# => romdata <= X"C407BFB4";
    when 16#0E13# => romdata <= X"82008001";
    when 16#0E14# => romdata <= X"C227BFB4";
    when 16#0E15# => romdata <= X"C207BFB0";
    when 16#0E16# => romdata <= X"82006001";
    when 16#0E17# => romdata <= X"C227BFB0";
    when 16#0E18# => romdata <= X"80A06007";
    when 16#0E19# => romdata <= X"04BFFEB8";
    when 16#0E1A# => romdata <= X"A0042008";
    when 16#0E1B# => romdata <= X"90100019";
    when 16#0E1C# => romdata <= X"7FFFFE38";
    when 16#0E1D# => romdata <= X"9207BFAC";
    when 16#0E1E# => romdata <= X"80A22000";
    when 16#0E1F# => romdata <= X"128000B2";
    when 16#0E20# => romdata <= X"C24FBFFF";
    when 16#0E21# => romdata <= X"80A06000";
    when 16#0E22# => romdata <= X"12BFFEB3";
    when 16#0E23# => romdata <= X"A0100013";
    when 16#0E24# => romdata <= X"808D2002";
    when 16#0E25# => romdata <= X"02BFFEBE";
    when 16#0E26# => romdata <= X"C207B90C";
    when 16#0E27# => romdata <= X"EA2FBFF9";
    when 16#0E28# => romdata <= X"82102030";
    when 16#0E29# => romdata <= X"C22FBFF8";
    when 16#0E2A# => romdata <= X"82102002";
    when 16#0E2B# => romdata <= X"C2242004";
    when 16#0E2C# => romdata <= X"8207BFF8";
    when 16#0E2D# => romdata <= X"C2240000";
    when 16#0E2E# => romdata <= X"C407BFB4";
    when 16#0E2F# => romdata <= X"C207BFB0";
    when 16#0E30# => romdata <= X"82006001";
    when 16#0E31# => romdata <= X"8400A002";
    when 16#0E32# => romdata <= X"C227BFB0";
    when 16#0E33# => romdata <= X"C427BFB4";
    when 16#0E34# => romdata <= X"80A06007";
    when 16#0E35# => romdata <= X"04BFFEAD";
    when 16#0E36# => romdata <= X"A0042008";
    when 16#0E37# => romdata <= X"90100019";
    when 16#0E38# => romdata <= X"7FFFFE1C";
    when 16#0E39# => romdata <= X"9207BFAC";
    when 16#0E3A# => romdata <= X"80A22000";
    when 16#0E3B# => romdata <= X"12800096";
    when 16#0E3C# => romdata <= X"C207B90C";
    when 16#0E3D# => romdata <= X"80A06080";
    when 16#0E3E# => romdata <= X"12BFFEA8";
    when 16#0E3F# => romdata <= X"A0100013";
    when 16#0E40# => romdata <= X"C407B910";
    when 16#0E41# => romdata <= X"82270002";
    when 16#0E42# => romdata <= X"80A06000";
    when 16#0E43# => romdata <= X"04BFFEA3";
    when 16#0E44# => romdata <= X"80A06010";
    when 16#0E45# => romdata <= X"04800024";
    when 16#0E46# => romdata <= X"E227B90C";
    when 16#0E47# => romdata <= X"86100010";
    when 16#0E48# => romdata <= X"84102010";
    when 16#0E49# => romdata <= X"A0100001";
    when 16#0E4A# => romdata <= X"10800006";
    when 16#0E4B# => romdata <= X"82100003";
    when 16#0E4C# => romdata <= X"A0043FF0";
    when 16#0E4D# => romdata <= X"80A42010";
    when 16#0E4E# => romdata <= X"24800019";
    when 16#0E4F# => romdata <= X"84100001";
    when 16#0E50# => romdata <= X"C4206004";
    when 16#0E51# => romdata <= X"E2204000";
    when 16#0E52# => romdata <= X"82006008";
    when 16#0E53# => romdata <= X"C607BFB0";
    when 16#0E54# => romdata <= X"C807BFB4";
    when 16#0E55# => romdata <= X"8600E001";
    when 16#0E56# => romdata <= X"88012010";
    when 16#0E57# => romdata <= X"C627BFB0";
    when 16#0E58# => romdata <= X"80A0E007";
    when 16#0E59# => romdata <= X"04BFFFF3";
    when 16#0E5A# => romdata <= X"C827BFB4";
    when 16#0E5B# => romdata <= X"C427B8E4";
    when 16#0E5C# => romdata <= X"90100019";
    when 16#0E5D# => romdata <= X"7FFFFDF7";
    when 16#0E5E# => romdata <= X"9207BFAC";
    when 16#0E5F# => romdata <= X"80A22000";
    when 16#0E60# => romdata <= X"12800071";
    when 16#0E61# => romdata <= X"C407B8E4";
    when 16#0E62# => romdata <= X"A0043FF0";
    when 16#0E63# => romdata <= X"80A42010";
    when 16#0E64# => romdata <= X"14BFFFEC";
    when 16#0E65# => romdata <= X"82100013";
    when 16#0E66# => romdata <= X"84100001";
    when 16#0E67# => romdata <= X"82100010";
    when 16#0E68# => romdata <= X"A0100002";
    when 16#0E69# => romdata <= X"C2242004";
    when 16#0E6A# => romdata <= X"C607B90C";
    when 16#0E6B# => romdata <= X"C6240000";
    when 16#0E6C# => romdata <= X"C407BFB4";
    when 16#0E6D# => romdata <= X"82008001";
    when 16#0E6E# => romdata <= X"C227BFB4";
    when 16#0E6F# => romdata <= X"C207BFB0";
    when 16#0E70# => romdata <= X"82006001";
    when 16#0E71# => romdata <= X"C227BFB0";
    when 16#0E72# => romdata <= X"80A06007";
    when 16#0E73# => romdata <= X"04BFFE73";
    when 16#0E74# => romdata <= X"A0042008";
    when 16#0E75# => romdata <= X"90100019";
    when 16#0E76# => romdata <= X"7FFFFDDE";
    when 16#0E77# => romdata <= X"9207BFAC";
    when 16#0E78# => romdata <= X"80A22000";
    when 16#0E79# => romdata <= X"12800058";
    when 16#0E7A# => romdata <= X"A0100013";
    when 16#0E7B# => romdata <= X"10BFFE6C";
    when 16#0E7C# => romdata <= X"C407B908";
    when 16#0E7D# => romdata <= X"048000AC";
    when 16#0E7E# => romdata <= X"C207B8F4";
    when 16#0E7F# => romdata <= X"03100032";
    when 16#0E80# => romdata <= X"D51FB8F8";
    when 16#0E81# => romdata <= X"82106060";
    when 16#0E82# => romdata <= X"D1184000";
    when 16#0E83# => romdata <= X"81AA8A48";
    when 16#0E84# => romdata <= X"01000000";
    when 16#0E85# => romdata <= X"038000F8";
    when 16#0E86# => romdata <= X"C207BFF4";
    when 16#0E87# => romdata <= X"82102001";
    when 16#0E88# => romdata <= X"C2242004";
    when 16#0E89# => romdata <= X"03100032";
    when 16#0E8A# => romdata <= X"82106048";
    when 16#0E8B# => romdata <= X"C407BFB4";
    when 16#0E8C# => romdata <= X"C2240000";
    when 16#0E8D# => romdata <= X"C207BFB0";
    when 16#0E8E# => romdata <= X"82006001";
    when 16#0E8F# => romdata <= X"8400A001";
    when 16#0E90# => romdata <= X"C227BFB0";
    when 16#0E91# => romdata <= X"C427BFB4";
    when 16#0E92# => romdata <= X"80A06007";
    when 16#0E93# => romdata <= X"14800313";
    when 16#0E94# => romdata <= X"A0042008";
    when 16#0E95# => romdata <= X"C207BFF4";
    when 16#0E96# => romdata <= X"C407B8F4";
    when 16#0E97# => romdata <= X"80A04002";
    when 16#0E98# => romdata <= X"06800006";
    when 16#0E99# => romdata <= X"82102001";
    when 16#0E9A# => romdata <= X"808D2001";
    when 16#0E9B# => romdata <= X"02BFFE95";
    when 16#0E9C# => romdata <= X"808D2004";
    when 16#0E9D# => romdata <= X"82102001";
    when 16#0E9E# => romdata <= X"C2242004";
    when 16#0E9F# => romdata <= X"C607B8E8";
    when 16#0EA0# => romdata <= X"C6240000";
    when 16#0EA1# => romdata <= X"C207BFB0";
    when 16#0EA2# => romdata <= X"C407BFB4";
    when 16#0EA3# => romdata <= X"82006001";
    when 16#0EA4# => romdata <= X"8400A001";
    when 16#0EA5# => romdata <= X"C227BFB0";
    when 16#0EA6# => romdata <= X"C427BFB4";
    when 16#0EA7# => romdata <= X"80A06007";
    when 16#0EA8# => romdata <= X"14800406";
    when 16#0EA9# => romdata <= X"A0042008";
    when 16#0EAA# => romdata <= X"C207B8F4";
    when 16#0EAB# => romdata <= X"AA007FFF";
    when 16#0EAC# => romdata <= X"80A56000";
    when 16#0EAD# => romdata <= X"04BFFE82";
    when 16#0EAE# => romdata <= X"80A56010";
    when 16#0EAF# => romdata <= X"04800274";
    when 16#0EB0# => romdata <= X"E227B90C";
    when 16#0EB1# => romdata <= X"AE102010";
    when 16#0EB2# => romdata <= X"10800006";
    when 16#0EB3# => romdata <= X"BA07BFAC";
    when 16#0EB4# => romdata <= X"AA057FF0";
    when 16#0EB5# => romdata <= X"80A56010";
    when 16#0EB6# => romdata <= X"2480026E";
    when 16#0EB7# => romdata <= X"EA242004";
    when 16#0EB8# => romdata <= X"EE242004";
    when 16#0EB9# => romdata <= X"E2240000";
    when 16#0EBA# => romdata <= X"A0042008";
    when 16#0EBB# => romdata <= X"C207BFB0";
    when 16#0EBC# => romdata <= X"C407BFB4";
    when 16#0EBD# => romdata <= X"82006001";
    when 16#0EBE# => romdata <= X"8400A010";
    when 16#0EBF# => romdata <= X"C227BFB0";
    when 16#0EC0# => romdata <= X"80A06007";
    when 16#0EC1# => romdata <= X"04BFFFF3";
    when 16#0EC2# => romdata <= X"C427BFB4";
    when 16#0EC3# => romdata <= X"90100019";
    when 16#0EC4# => romdata <= X"7FFFFD90";
    when 16#0EC5# => romdata <= X"9210001D";
    when 16#0EC6# => romdata <= X"80A22000";
    when 16#0EC7# => romdata <= X"1280000A";
    when 16#0EC8# => romdata <= X"A0100013";
    when 16#0EC9# => romdata <= X"10BFFFEC";
    when 16#0ECA# => romdata <= X"AA057FF0";
    when 16#0ECB# => romdata <= X"90100019";
    when 16#0ECC# => romdata <= X"7FFFFD88";
    when 16#0ECD# => romdata <= X"9207BFAC";
    when 16#0ECE# => romdata <= X"80A22000";
    when 16#0ECF# => romdata <= X"22BFFE9F";
    when 16#0ED0# => romdata <= X"C027BFB0";
    when 16#0ED1# => romdata <= X"80A5A000";
    when 16#0ED2# => romdata <= X"22800006";
    when 16#0ED3# => romdata <= X"C216600C";
    when 16#0ED4# => romdata <= X"D007A044";
    when 16#0ED5# => romdata <= X"40000D62";
    when 16#0ED6# => romdata <= X"92100016";
    when 16#0ED7# => romdata <= X"C216600C";
    when 16#0ED8# => romdata <= X"83286010";
    when 16#0ED9# => romdata <= X"83306010";
    when 16#0EDA# => romdata <= X"80886200";
    when 16#0EDB# => romdata <= X"0280009E";
    when 16#0EDC# => romdata <= X"01000000";
    when 16#0EDD# => romdata <= X"80886040";
    when 16#0EDE# => romdata <= X"12800004";
    when 16#0EDF# => romdata <= X"01000000";
    when 16#0EE0# => romdata <= X"81C7E008";
    when 16#0EE1# => romdata <= X"81E80000";
    when 16#0EE2# => romdata <= X"81C7E008";
    when 16#0EE3# => romdata <= X"91E83FFF";
    when 16#0EE4# => romdata <= X"40000659";
    when 16#0EE5# => romdata <= X"90100019";
    when 16#0EE6# => romdata <= X"80A22000";
    when 16#0EE7# => romdata <= X"3280041D";
    when 16#0EE8# => romdata <= X"C216600C";
    when 16#0EE9# => romdata <= X"C616600C";
    when 16#0EEA# => romdata <= X"82100003";
    when 16#0EEB# => romdata <= X"8408E01A";
    when 16#0EEC# => romdata <= X"80A0A00A";
    when 16#0EED# => romdata <= X"12BFFD93";
    when 16#0EEE# => romdata <= X"A607BF40";
    when 16#0EEF# => romdata <= X"C456600E";
    when 16#0EF0# => romdata <= X"80A0A000";
    when 16#0EF1# => romdata <= X"06BFFD8E";
    when 16#0EF2# => romdata <= X"C416600E";
    when 16#0EF3# => romdata <= X"80886200";
    when 16#0EF4# => romdata <= X"028000E6";
    when 16#0EF5# => romdata <= X"01000000";
    when 16#0EF6# => romdata <= X"8608FFFD";
    when 16#0EF7# => romdata <= X"C2066024";
    when 16#0EF8# => romdata <= X"C227BE98";
    when 16#0EF9# => romdata <= X"8207B918";
    when 16#0EFA# => romdata <= X"C806601C";
    when 16#0EFB# => romdata <= X"C227BE84";
    when 16#0EFC# => romdata <= X"C227BE74";
    when 16#0EFD# => romdata <= X"82102400";
    when 16#0EFE# => romdata <= X"C637BE80";
    when 16#0EFF# => romdata <= X"C437BE82";
    when 16#0F00# => romdata <= X"C827BE90";
    when 16#0F01# => romdata <= X"A207BF80";
    when 16#0F02# => romdata <= X"C227BE88";
    when 16#0F03# => romdata <= X"C227BE7C";
    when 16#0F04# => romdata <= X"90100011";
    when 16#0F05# => romdata <= X"40001BC0";
    when 16#0F06# => romdata <= X"C027BE8C";
    when 16#0F07# => romdata <= X"90100011";
    when 16#0F08# => romdata <= X"40001BD3";
    when 16#0F09# => romdata <= X"92102001";
    when 16#0F0A# => romdata <= X"92100011";
    when 16#0F0B# => romdata <= X"A007BECC";
    when 16#0F0C# => romdata <= X"40001B80";
    when 16#0F0D# => romdata <= X"90100010";
    when 16#0F0E# => romdata <= X"40001BC2";
    when 16#0F0F# => romdata <= X"90100011";
    when 16#0F10# => romdata <= X"D007A044";
    when 16#0F11# => romdata <= X"A207BE74";
    when 16#0F12# => romdata <= X"9410001A";
    when 16#0F13# => romdata <= X"92100011";
    when 16#0F14# => romdata <= X"7FFFFD4E";
    when 16#0F15# => romdata <= X"9610001B";
    when 16#0F16# => romdata <= X"B0922000";
    when 16#0F17# => romdata <= X"06800008";
    when 16#0F18# => romdata <= X"C217BE80";
    when 16#0F19# => romdata <= X"40000BB8";
    when 16#0F1A# => romdata <= X"90100011";
    when 16#0F1B# => romdata <= X"80A22000";
    when 16#0F1C# => romdata <= X"32800002";
    when 16#0F1D# => romdata <= X"B0103FFF";
    when 16#0F1E# => romdata <= X"C217BE80";
    when 16#0F1F# => romdata <= X"80886040";
    when 16#0F20# => romdata <= X"02800005";
    when 16#0F21# => romdata <= X"01000000";
    when 16#0F22# => romdata <= X"C216600C";
    when 16#0F23# => romdata <= X"82106040";
    when 16#0F24# => romdata <= X"C236600C";
    when 16#0F25# => romdata <= X"40001B74";
    when 16#0F26# => romdata <= X"90100010";
    when 16#0F27# => romdata <= X"81C7E008";
    when 16#0F28# => romdata <= X"81E80000";
    when 16#0F29# => romdata <= X"80A06001";
    when 16#0F2A# => romdata <= X"048001B6";
    when 16#0F2B# => romdata <= X"808D2001";
    when 16#0F2C# => romdata <= X"C20DC000";
    when 16#0F2D# => romdata <= X"C22FBFF8";
    when 16#0F2E# => romdata <= X"8210202E";
    when 16#0F2F# => romdata <= X"C22FBFF9";
    when 16#0F30# => romdata <= X"82102002";
    when 16#0F31# => romdata <= X"C2242004";
    when 16#0F32# => romdata <= X"8207BFF8";
    when 16#0F33# => romdata <= X"C2240000";
    when 16#0F34# => romdata <= X"C407BFB4";
    when 16#0F35# => romdata <= X"C207BFB0";
    when 16#0F36# => romdata <= X"82006001";
    when 16#0F37# => romdata <= X"8400A002";
    when 16#0F38# => romdata <= X"C227BFB0";
    when 16#0F39# => romdata <= X"C427BFB4";
    when 16#0F3A# => romdata <= X"80A06007";
    when 16#0F3B# => romdata <= X"148001BB";
    when 16#0F3C# => romdata <= X"A0042008";
    when 16#0F3D# => romdata <= X"05100032";
    when 16#0F3E# => romdata <= X"D51FB8F8";
    when 16#0F3F# => romdata <= X"8410A060";
    when 16#0F40# => romdata <= X"D1188000";
    when 16#0F41# => romdata <= X"81AA8A48";
    when 16#0F42# => romdata <= X"01000000";
    when 16#0F43# => romdata <= X"13800072";
    when 16#0F44# => romdata <= X"C607B8F4";
    when 16#0F45# => romdata <= X"C407B8F4";
    when 16#0F46# => romdata <= X"8200BFFF";
    when 16#0F47# => romdata <= X"C2242004";
    when 16#0F48# => romdata <= X"AE05E001";
    when 16#0F49# => romdata <= X"EE240000";
    when 16#0F4A# => romdata <= X"C407BFB4";
    when 16#0F4B# => romdata <= X"82008001";
    when 16#0F4C# => romdata <= X"C227BFB4";
    when 16#0F4D# => romdata <= X"C207BFB0";
    when 16#0F4E# => romdata <= X"82006001";
    when 16#0F4F# => romdata <= X"C227BFB0";
    when 16#0F50# => romdata <= X"80A06007";
    when 16#0F51# => romdata <= X"1480019D";
    when 16#0F52# => romdata <= X"A0042008";
    when 16#0F53# => romdata <= X"C407B8F0";
    when 16#0F54# => romdata <= X"C4242004";
    when 16#0F55# => romdata <= X"8207BFE0";
    when 16#0F56# => romdata <= X"C607B8F0";
    when 16#0F57# => romdata <= X"C2240000";
    when 16#0F58# => romdata <= X"C407BFB4";
    when 16#0F59# => romdata <= X"C207BFB0";
    when 16#0F5A# => romdata <= X"82006001";
    when 16#0F5B# => romdata <= X"84008003";
    when 16#0F5C# => romdata <= X"C427BFB4";
    when 16#0F5D# => romdata <= X"C227BFB0";
    when 16#0F5E# => romdata <= X"80A06007";
    when 16#0F5F# => romdata <= X"04BFFDD0";
    when 16#0F60# => romdata <= X"A0042008";
    when 16#0F61# => romdata <= X"90100019";
    when 16#0F62# => romdata <= X"7FFFFCF2";
    when 16#0F63# => romdata <= X"9207BFAC";
    when 16#0F64# => romdata <= X"80A22000";
    when 16#0F65# => romdata <= X"12BFFF6C";
    when 16#0F66# => romdata <= X"A0100013";
    when 16#0F67# => romdata <= X"10BFFDC9";
    when 16#0F68# => romdata <= X"808D2004";
    when 16#0F69# => romdata <= X"90100019";
    when 16#0F6A# => romdata <= X"7FFFFCEA";
    when 16#0F6B# => romdata <= X"9207BFAC";
    when 16#0F6C# => romdata <= X"80A22000";
    when 16#0F6D# => romdata <= X"12BFFF6A";
    when 16#0F6E# => romdata <= X"A0100013";
    when 16#0F6F# => romdata <= X"10BFFD3C";
    when 16#0F70# => romdata <= X"C20D0000";
    when 16#0F71# => romdata <= X"40001B33";
    when 16#0F72# => romdata <= X"90066058";
    when 16#0F73# => romdata <= X"10BFFCF9";
    when 16#0F74# => romdata <= X"03100032";
    when 16#0F75# => romdata <= X"40000C11";
    when 16#0F76# => romdata <= X"01000000";
    when 16#0F77# => romdata <= X"10BFFCFE";
    when 16#0F78# => romdata <= X"C216600C";
    when 16#0F79# => romdata <= X"40001B41";
    when 16#0F7A# => romdata <= X"90066058";
    when 16#0F7B# => romdata <= X"10BFFF62";
    when 16#0F7C# => romdata <= X"C216600C";
    when 16#0F7D# => romdata <= X"80A06000";
    when 16#0F7E# => romdata <= X"04800239";
    when 16#0F7F# => romdata <= X"C407B8F4";
    when 16#0F80# => romdata <= X"80A04002";
    when 16#0F81# => romdata <= X"268001DD";
    when 16#0F82# => romdata <= X"C2242004";
    when 16#0F83# => romdata <= X"C4242004";
    when 16#0F84# => romdata <= X"C607B8F4";
    when 16#0F85# => romdata <= X"EE240000";
    when 16#0F86# => romdata <= X"C207BFB0";
    when 16#0F87# => romdata <= X"C407BFB4";
    when 16#0F88# => romdata <= X"82006001";
    when 16#0F89# => romdata <= X"84008003";
    when 16#0F8A# => romdata <= X"C227BFB0";
    when 16#0F8B# => romdata <= X"C427BFB4";
    when 16#0F8C# => romdata <= X"80A06007";
    when 16#0F8D# => romdata <= X"1480026F";
    when 16#0F8E# => romdata <= X"A0042008";
    when 16#0F8F# => romdata <= X"EA07BFF4";
    when 16#0F90# => romdata <= X"C207B8F4";
    when 16#0F91# => romdata <= X"AA254001";
    when 16#0F92# => romdata <= X"80A56000";
    when 16#0F93# => romdata <= X"04800201";
    when 16#0F94# => romdata <= X"80A56010";
    when 16#0F95# => romdata <= X"048001ED";
    when 16#0F96# => romdata <= X"E227B90C";
    when 16#0F97# => romdata <= X"AE102010";
    when 16#0F98# => romdata <= X"10800006";
    when 16#0F99# => romdata <= X"BA07BFAC";
    when 16#0F9A# => romdata <= X"AA057FF0";
    when 16#0F9B# => romdata <= X"80A56010";
    when 16#0F9C# => romdata <= X"248001E7";
    when 16#0F9D# => romdata <= X"EA242004";
    when 16#0F9E# => romdata <= X"EE242004";
    when 16#0F9F# => romdata <= X"E2240000";
    when 16#0FA0# => romdata <= X"A0042008";
    when 16#0FA1# => romdata <= X"C207BFB0";
    when 16#0FA2# => romdata <= X"C407BFB4";
    when 16#0FA3# => romdata <= X"82006001";
    when 16#0FA4# => romdata <= X"8400A010";
    when 16#0FA5# => romdata <= X"C227BFB0";
    when 16#0FA6# => romdata <= X"80A06007";
    when 16#0FA7# => romdata <= X"04BFFFF3";
    when 16#0FA8# => romdata <= X"C427BFB4";
    when 16#0FA9# => romdata <= X"90100019";
    when 16#0FAA# => romdata <= X"7FFFFCAA";
    when 16#0FAB# => romdata <= X"9210001D";
    when 16#0FAC# => romdata <= X"80A22000";
    when 16#0FAD# => romdata <= X"12BFFF24";
    when 16#0FAE# => romdata <= X"A0100013";
    when 16#0FAF# => romdata <= X"10BFFFEC";
    when 16#0FB0# => romdata <= X"AA057FF0";
    when 16#0FB1# => romdata <= X"AE07BE73";
    when 16#0FB2# => romdata <= X"C22FBE73";
    when 16#0FB3# => romdata <= X"10BFFE23";
    when 16#0FB4# => romdata <= X"BA102001";
    when 16#0FB5# => romdata <= X"AA00FFFF";
    when 16#0FB6# => romdata <= X"80A56000";
    when 16#0FB7# => romdata <= X"04BFFF9C";
    when 16#0FB8# => romdata <= X"80A56010";
    when 16#0FB9# => romdata <= X"04800145";
    when 16#0FBA# => romdata <= X"E227B90C";
    when 16#0FBB# => romdata <= X"AE102010";
    when 16#0FBC# => romdata <= X"10800006";
    when 16#0FBD# => romdata <= X"BA07BFAC";
    when 16#0FBE# => romdata <= X"AA057FF0";
    when 16#0FBF# => romdata <= X"80A56010";
    when 16#0FC0# => romdata <= X"2480013F";
    when 16#0FC1# => romdata <= X"EA242004";
    when 16#0FC2# => romdata <= X"EE242004";
    when 16#0FC3# => romdata <= X"E2240000";
    when 16#0FC4# => romdata <= X"A0042008";
    when 16#0FC5# => romdata <= X"C207BFB0";
    when 16#0FC6# => romdata <= X"C407BFB4";
    when 16#0FC7# => romdata <= X"82006001";
    when 16#0FC8# => romdata <= X"8400A010";
    when 16#0FC9# => romdata <= X"C227BFB0";
    when 16#0FCA# => romdata <= X"80A06007";
    when 16#0FCB# => romdata <= X"04BFFFF3";
    when 16#0FCC# => romdata <= X"C427BFB4";
    when 16#0FCD# => romdata <= X"90100019";
    when 16#0FCE# => romdata <= X"7FFFFC86";
    when 16#0FCF# => romdata <= X"9210001D";
    when 16#0FD0# => romdata <= X"80A22000";
    when 16#0FD1# => romdata <= X"12BFFF00";
    when 16#0FD2# => romdata <= X"A0100013";
    when 16#0FD3# => romdata <= X"10BFFFEC";
    when 16#0FD4# => romdata <= X"AA057FF0";
    when 16#0FD5# => romdata <= X"22BFFDF3";
    when 16#0FD6# => romdata <= X"FA06C000";
    when 16#0FD7# => romdata <= X"FA56E002";
    when 16#0FD8# => romdata <= X"10BFFDF1";
    when 16#0FD9# => romdata <= X"B606E004";
    when 16#0FDA# => romdata <= X"40001AE0";
    when 16#0FDB# => romdata <= X"90066058";
    when 16#0FDC# => romdata <= X"C616600C";
    when 16#0FDD# => romdata <= X"10BFFF19";
    when 16#0FDE# => romdata <= X"C416600E";
    when 16#0FDF# => romdata <= X"F806C000";
    when 16#0FE0# => romdata <= X"80A72000";
    when 16#0FE1# => romdata <= X"16800026";
    when 16#0FE2# => romdata <= X"B606E004";
    when 16#0FE3# => romdata <= X"B820001C";
    when 16#0FE4# => romdata <= X"EA0E8000";
    when 16#0FE5# => romdata <= X"A8152004";
    when 16#0FE6# => romdata <= X"10BFFCD3";
    when 16#0FE7# => romdata <= X"AB2D6018";
    when 16#0FE8# => romdata <= X"80A56043";
    when 16#0FE9# => romdata <= X"02800123";
    when 16#0FEA# => romdata <= X"808D2010";
    when 16#0FEB# => romdata <= X"32800122";
    when 16#0FEC# => romdata <= X"AC07BFD8";
    when 16#0FED# => romdata <= X"C206C000";
    when 16#0FEE# => romdata <= X"BA102001";
    when 16#0FEF# => romdata <= X"B606E004";
    when 16#0FF0# => romdata <= X"AE07BD18";
    when 16#0FF1# => romdata <= X"C22FBD18";
    when 16#0FF2# => romdata <= X"8238001D";
    when 16#0FF3# => romdata <= X"C02FBFFF";
    when 16#0FF4# => romdata <= X"8338601F";
    when 16#0FF5# => romdata <= X"C027B908";
    when 16#0FF6# => romdata <= X"820F4001";
    when 16#0FF7# => romdata <= X"AC102000";
    when 16#0FF8# => romdata <= X"10BFFCD1";
    when 16#0FF9# => romdata <= X"C227B910";
    when 16#0FFA# => romdata <= X"808D2010";
    when 16#0FFB# => romdata <= X"128000C0";
    when 16#0FFC# => romdata <= X"C206C000";
    when 16#0FFD# => romdata <= X"808D2040";
    when 16#0FFE# => romdata <= X"028000BD";
    when 16#0FFF# => romdata <= X"01000000";
    when 16#1000# => romdata <= X"B606E004";
    when 16#1001# => romdata <= X"10BFFC8C";
    when 16#1002# => romdata <= X"F0304000";
    when 16#1003# => romdata <= X"EA0E8000";
    when 16#1004# => romdata <= X"A8152001";
    when 16#1005# => romdata <= X"10BFFCB4";
    when 16#1006# => romdata <= X"AB2D6018";
    when 16#1007# => romdata <= X"EA0E8000";
    when 16#1008# => romdata <= X"10BFFCB1";
    when 16#1009# => romdata <= X"AB2D6018";
    when 16#100A# => romdata <= X"C62FBFFF";
    when 16#100B# => romdata <= X"EA0E8000";
    when 16#100C# => romdata <= X"10BFFCAD";
    when 16#100D# => romdata <= X"AB2D6018";
    when 16#100E# => romdata <= X"EA0E8000";
    when 16#100F# => romdata <= X"A8152080";
    when 16#1010# => romdata <= X"10BFFCA9";
    when 16#1011# => romdata <= X"AB2D6018";
    when 16#1012# => romdata <= X"82057FD0";
    when 16#1013# => romdata <= X"B8102000";
    when 16#1014# => romdata <= X"EA4E8000";
    when 16#1015# => romdata <= X"852F2003";
    when 16#1016# => romdata <= X"B92F2001";
    when 16#1017# => romdata <= X"B8070002";
    when 16#1018# => romdata <= X"B800401C";
    when 16#1019# => romdata <= X"82057FD0";
    when 16#101A# => romdata <= X"80A06009";
    when 16#101B# => romdata <= X"08BFFFF9";
    when 16#101C# => romdata <= X"B406A001";
    when 16#101D# => romdata <= X"10BFFC9F";
    when 16#101E# => romdata <= X"82057FE0";
    when 16#101F# => romdata <= X"FA06C000";
    when 16#1020# => romdata <= X"80A0001D";
    when 16#1021# => romdata <= X"07100032";
    when 16#1022# => romdata <= X"B606E004";
    when 16#1023# => romdata <= X"8610E028";
    when 16#1024# => romdata <= X"84402000";
    when 16#1025# => romdata <= X"A8152002";
    when 16#1026# => romdata <= X"C627B8EC";
    when 16#1027# => romdata <= X"82102002";
    when 16#1028# => romdata <= X"10BFFD61";
    when 16#1029# => romdata <= X"AA102078";
    when 16#102A# => romdata <= X"EA0E8000";
    when 16#102B# => romdata <= X"A8152010";
    when 16#102C# => romdata <= X"10BFFC8D";
    when 16#102D# => romdata <= X"AB2D6018";
    when 16#102E# => romdata <= X"EA0E8000";
    when 16#102F# => romdata <= X"AB2D6018";
    when 16#1030# => romdata <= X"833D6018";
    when 16#1031# => romdata <= X"80A0606C";
    when 16#1032# => romdata <= X"22800204";
    when 16#1033# => romdata <= X"B406A001";
    when 16#1034# => romdata <= X"10BFFC85";
    when 16#1035# => romdata <= X"A8152010";
    when 16#1036# => romdata <= X"03100032";
    when 16#1037# => romdata <= X"82106028";
    when 16#1038# => romdata <= X"808D2010";
    when 16#1039# => romdata <= X"1280004E";
    when 16#103A# => romdata <= X"C227B8EC";
    when 16#103B# => romdata <= X"808D2040";
    when 16#103C# => romdata <= X"2280004C";
    when 16#103D# => romdata <= X"FA06C000";
    when 16#103E# => romdata <= X"FA16E002";
    when 16#103F# => romdata <= X"B606E004";
    when 16#1040# => romdata <= X"80A0001D";
    when 16#1041# => romdata <= X"84402000";
    when 16#1042# => romdata <= X"80A0A000";
    when 16#1043# => romdata <= X"02BFFD46";
    when 16#1044# => romdata <= X"82102002";
    when 16#1045# => romdata <= X"808D2001";
    when 16#1046# => romdata <= X"22BFFD44";
    when 16#1047# => romdata <= X"C02FBFFF";
    when 16#1048# => romdata <= X"A8152002";
    when 16#1049# => romdata <= X"10BFFD40";
    when 16#104A# => romdata <= X"84102001";
    when 16#104B# => romdata <= X"EA4E8000";
    when 16#104C# => romdata <= X"80A5602A";
    when 16#104D# => romdata <= X"02800348";
    when 16#104E# => romdata <= X"B406A001";
    when 16#104F# => romdata <= X"82057FD0";
    when 16#1050# => romdata <= X"84102000";
    when 16#1051# => romdata <= X"80A06009";
    when 16#1052# => romdata <= X"18BFFC69";
    when 16#1053# => romdata <= X"AC102000";
    when 16#1054# => romdata <= X"EA4E8000";
    when 16#1055# => romdata <= X"9B28A003";
    when 16#1056# => romdata <= X"8528A001";
    when 16#1057# => romdata <= X"8400800D";
    when 16#1058# => romdata <= X"84008001";
    when 16#1059# => romdata <= X"82057FD0";
    when 16#105A# => romdata <= X"80A06009";
    when 16#105B# => romdata <= X"08BFFFF9";
    when 16#105C# => romdata <= X"B406A001";
    when 16#105D# => romdata <= X"AC90A000";
    when 16#105E# => romdata <= X"26BFFC5D";
    when 16#105F# => romdata <= X"AC103FFF";
    when 16#1060# => romdata <= X"10BFFC5C";
    when 16#1061# => romdata <= X"82057FE0";
    when 16#1062# => romdata <= X"EA0E8000";
    when 16#1063# => romdata <= X"A8152040";
    when 16#1064# => romdata <= X"10BFFC55";
    when 16#1065# => romdata <= X"AB2D6018";
    when 16#1066# => romdata <= X"C02FBFFF";
    when 16#1067# => romdata <= X"EE06C000";
    when 16#1068# => romdata <= X"80A5E000";
    when 16#1069# => romdata <= X"02800273";
    when 16#106A# => romdata <= X"B606E004";
    when 16#106B# => romdata <= X"80A56053";
    when 16#106C# => romdata <= X"028000C7";
    when 16#106D# => romdata <= X"808D2010";
    when 16#106E# => romdata <= X"328000C6";
    when 16#106F# => romdata <= X"EE27BFF0";
    when 16#1070# => romdata <= X"80A5A000";
    when 16#1071# => romdata <= X"068001AB";
    when 16#1072# => romdata <= X"90100017";
    when 16#1073# => romdata <= X"92102000";
    when 16#1074# => romdata <= X"40000E67";
    when 16#1075# => romdata <= X"94100016";
    when 16#1076# => romdata <= X"80A22000";
    when 16#1077# => romdata <= X"22800007";
    when 16#1078# => romdata <= X"EC27B910";
    when 16#1079# => romdata <= X"BA220017";
    when 16#107A# => romdata <= X"80A74016";
    when 16#107B# => romdata <= X"0480023B";
    when 16#107C# => romdata <= X"8238001D";
    when 16#107D# => romdata <= X"EC27B910";
    when 16#107E# => romdata <= X"BA100016";
    when 16#107F# => romdata <= X"C027B908";
    when 16#1080# => romdata <= X"10BFFD5C";
    when 16#1081# => romdata <= X"AC102000";
    when 16#1082# => romdata <= X"07100032";
    when 16#1083# => romdata <= X"8610E008";
    when 16#1084# => romdata <= X"808D2010";
    when 16#1085# => romdata <= X"02BFFFB6";
    when 16#1086# => romdata <= X"C627B8EC";
    when 16#1087# => romdata <= X"FA06C000";
    when 16#1088# => romdata <= X"10BFFFB8";
    when 16#1089# => romdata <= X"B606E004";
    when 16#108A# => romdata <= X"C24FBFFF";
    when 16#108B# => romdata <= X"80A06000";
    when 16#108C# => romdata <= X"32BFFF7C";
    when 16#108D# => romdata <= X"EA0E8000";
    when 16#108E# => romdata <= X"C82FBFFF";
    when 16#108F# => romdata <= X"EA0E8000";
    when 16#1090# => romdata <= X"10BFFC29";
    when 16#1091# => romdata <= X"AB2D6018";
    when 16#1092# => romdata <= X"EA0E8000";
    when 16#1093# => romdata <= X"A8152008";
    when 16#1094# => romdata <= X"10BFFC25";
    when 16#1095# => romdata <= X"AB2D6018";
    when 16#1096# => romdata <= X"80A5BFFF";
    when 16#1097# => romdata <= X"0280019D";
    when 16#1098# => romdata <= X"80A56047";
    when 16#1099# => romdata <= X"02800108";
    when 16#109A# => romdata <= X"80A56067";
    when 16#109B# => romdata <= X"02800107";
    when 16#109C# => romdata <= X"80A5A000";
    when 16#109D# => romdata <= X"808D2008";
    when 16#109E# => romdata <= X"0280008D";
    when 16#109F# => romdata <= X"9210001B";
    when 16#10A0# => romdata <= X"9007BFC8";
    when 16#10A1# => romdata <= X"40000E76";
    when 16#10A2# => romdata <= X"94102008";
    when 16#10A3# => romdata <= X"D11FBFC8";
    when 16#10A4# => romdata <= X"D13FB8F8";
    when 16#10A5# => romdata <= X"D13FB910";
    when 16#10A6# => romdata <= X"B606E008";
    when 16#10A7# => romdata <= X"40001482";
    when 16#10A8# => romdata <= X"D01FB8F8";
    when 16#10A9# => romdata <= X"80A22000";
    when 16#10AA# => romdata <= X"02800190";
    when 16#10AB# => romdata <= X"03100032";
    when 16#10AC# => romdata <= X"D51FB8F8";
    when 16#10AD# => romdata <= X"82106060";
    when 16#10AE# => romdata <= X"D1184000";
    when 16#10AF# => romdata <= X"81AA8AC8";
    when 16#10B0# => romdata <= X"01000000";
    when 16#10B1# => romdata <= X"098000FD";
    when 16#10B2# => romdata <= X"8210202D";
    when 16#10B3# => romdata <= X"82102003";
    when 16#10B4# => romdata <= X"2F100032";
    when 16#10B5# => romdata <= X"C227B910";
    when 16#10B6# => romdata <= X"BA102003";
    when 16#10B7# => romdata <= X"C027B908";
    when 16#10B8# => romdata <= X"AE15E020";
    when 16#10B9# => romdata <= X"10BFFD23";
    when 16#10BA# => romdata <= X"AC102000";
    when 16#10BB# => romdata <= X"B606E004";
    when 16#10BC# => romdata <= X"10BFFBD1";
    when 16#10BD# => romdata <= X"F0204000";
    when 16#10BE# => romdata <= X"C407B8EC";
    when 16#10BF# => romdata <= X"820F600F";
    when 16#10C0# => romdata <= X"C2088001";
    when 16#10C1# => romdata <= X"AE05FFFF";
    when 16#10C2# => romdata <= X"BB376004";
    when 16#10C3# => romdata <= X"80A76000";
    when 16#10C4# => romdata <= X"12BFFFFB";
    when 16#10C5# => romdata <= X"C22DC000";
    when 16#10C6# => romdata <= X"C207B8DC";
    when 16#10C7# => romdata <= X"10BFFD0F";
    when 16#10C8# => romdata <= X"BA204017";
    when 16#10C9# => romdata <= X"80A76009";
    when 16#10CA# => romdata <= X"08800010";
    when 16#10CB# => romdata <= X"8407BE74";
    when 16#10CC# => romdata <= X"AE100002";
    when 16#10CD# => romdata <= X"9010001D";
    when 16#10CE# => romdata <= X"9210200A";
    when 16#10CF# => romdata <= X"400016A5";
    when 16#10D0# => romdata <= X"AE05FFFF";
    when 16#10D1# => romdata <= X"82022030";
    when 16#10D2# => romdata <= X"9210200A";
    when 16#10D3# => romdata <= X"9010001D";
    when 16#10D4# => romdata <= X"400015F4";
    when 16#10D5# => romdata <= X"C22DC000";
    when 16#10D6# => romdata <= X"80A22009";
    when 16#10D7# => romdata <= X"18BFFFF6";
    when 16#10D8# => romdata <= X"BA100008";
    when 16#10D9# => romdata <= X"84100017";
    when 16#10DA# => romdata <= X"82076030";
    when 16#10DB# => romdata <= X"C607B8DC";
    when 16#10DC# => romdata <= X"AE00BFFF";
    when 16#10DD# => romdata <= X"C228BFFF";
    when 16#10DE# => romdata <= X"10BFFCF8";
    when 16#10DF# => romdata <= X"BA20C017";
    when 16#10E0# => romdata <= X"32BFFE4D";
    when 16#10E1# => romdata <= X"C20DC000";
    when 16#10E2# => romdata <= X"82102001";
    when 16#10E3# => romdata <= X"C2242004";
    when 16#10E4# => romdata <= X"EE240000";
    when 16#10E5# => romdata <= X"A0042008";
    when 16#10E6# => romdata <= X"C207BFB0";
    when 16#10E7# => romdata <= X"C407BFB4";
    when 16#10E8# => romdata <= X"82006001";
    when 16#10E9# => romdata <= X"8400A001";
    when 16#10EA# => romdata <= X"C227BFB0";
    when 16#10EB# => romdata <= X"80A06007";
    when 16#10EC# => romdata <= X"04BFFE67";
    when 16#10ED# => romdata <= X"C427BFB4";
    when 16#10EE# => romdata <= X"90100019";
    when 16#10EF# => romdata <= X"7FFFFB65";
    when 16#10F0# => romdata <= X"9207BFAC";
    when 16#10F1# => romdata <= X"80A22000";
    when 16#10F2# => romdata <= X"12BFFDDF";
    when 16#10F3# => romdata <= X"A0100013";
    when 16#10F4# => romdata <= X"10BFFE60";
    when 16#10F5# => romdata <= X"C407B8F0";
    when 16#10F6# => romdata <= X"90100019";
    when 16#10F7# => romdata <= X"7FFFFB5D";
    when 16#10F8# => romdata <= X"9207BFAC";
    when 16#10F9# => romdata <= X"80A22000";
    when 16#10FA# => romdata <= X"12BFFDD7";
    when 16#10FB# => romdata <= X"A0100013";
    when 16#10FC# => romdata <= X"10BFFE42";
    when 16#10FD# => romdata <= X"05100032";
    when 16#10FE# => romdata <= X"EA242004";
    when 16#10FF# => romdata <= X"C207B90C";
    when 16#1100# => romdata <= X"C2240000";
    when 16#1101# => romdata <= X"C207BFB4";
    when 16#1102# => romdata <= X"AA004015";
    when 16#1103# => romdata <= X"C207BFB0";
    when 16#1104# => romdata <= X"82006001";
    when 16#1105# => romdata <= X"EA27BFB4";
    when 16#1106# => romdata <= X"C227BFB0";
    when 16#1107# => romdata <= X"80A06007";
    when 16#1108# => romdata <= X"04BFFE4B";
    when 16#1109# => romdata <= X"A0042008";
    when 16#110A# => romdata <= X"10BFFFE5";
    when 16#110B# => romdata <= X"90100019";
    when 16#110C# => romdata <= X"AC07BFD8";
    when 16#110D# => romdata <= X"92102000";
    when 16#110E# => romdata <= X"94102008";
    when 16#110F# => romdata <= X"40000E9B";
    when 16#1110# => romdata <= X"90100016";
    when 16#1111# => romdata <= X"D406C000";
    when 16#1112# => romdata <= X"D007A044";
    when 16#1113# => romdata <= X"96100016";
    when 16#1114# => romdata <= X"AE07BD18";
    when 16#1115# => romdata <= X"400002AD";
    when 16#1116# => romdata <= X"92100017";
    when 16#1117# => romdata <= X"80A23FFF";
    when 16#1118# => romdata <= X"02800228";
    when 16#1119# => romdata <= X"BA100008";
    when 16#111A# => romdata <= X"10BFFED8";
    when 16#111B# => romdata <= X"B606E004";
    when 16#111C# => romdata <= X"8210202D";
    when 16#111D# => romdata <= X"BA20001D";
    when 16#111E# => romdata <= X"C22FBFFF";
    when 16#111F# => romdata <= X"80A0001D";
    when 16#1120# => romdata <= X"82102001";
    when 16#1121# => romdata <= X"10BFFC69";
    when 16#1122# => romdata <= X"84402000";
    when 16#1123# => romdata <= X"EA242004";
    when 16#1124# => romdata <= X"C407B90C";
    when 16#1125# => romdata <= X"C4240000";
    when 16#1126# => romdata <= X"C207BFB4";
    when 16#1127# => romdata <= X"AA004015";
    when 16#1128# => romdata <= X"A0042008";
    when 16#1129# => romdata <= X"10BFFC01";
    when 16#112A# => romdata <= X"EA27BFB4";
    when 16#112B# => romdata <= X"9007BFC0";
    when 16#112C# => romdata <= X"40000DEB";
    when 16#112D# => romdata <= X"94102008";
    when 16#112E# => romdata <= X"D51FBFC0";
    when 16#112F# => romdata <= X"D53FB8F8";
    when 16#1130# => romdata <= X"B606E008";
    when 16#1131# => romdata <= X"10BFFF76";
    when 16#1132# => romdata <= X"D53FB910";
    when 16#1133# => romdata <= X"EE27BFF0";
    when 16#1134# => romdata <= X"92102000";
    when 16#1135# => romdata <= X"9007BFD0";
    when 16#1136# => romdata <= X"40000E74";
    when 16#1137# => romdata <= X"94102008";
    when 16#1138# => romdata <= X"80A5A000";
    when 16#1139# => romdata <= X"068001F4";
    when 16#113A# => romdata <= X"BA102000";
    when 16#113B# => romdata <= X"82102000";
    when 16#113C# => romdata <= X"F627B910";
    when 16#113D# => romdata <= X"B6100015";
    when 16#113E# => romdata <= X"AA100010";
    when 16#113F# => romdata <= X"A010001D";
    when 16#1140# => romdata <= X"BA100016";
    when 16#1141# => romdata <= X"10800003";
    when 16#1142# => romdata <= X"AC100001";
    when 16#1143# => romdata <= X"A0100001";
    when 16#1144# => romdata <= X"C207BFF0";
    when 16#1145# => romdata <= X"D4004016";
    when 16#1146# => romdata <= X"80A2A000";
    when 16#1147# => romdata <= X"028001C4";
    when 16#1148# => romdata <= X"D007A044";
    when 16#1149# => romdata <= X"9207BD18";
    when 16#114A# => romdata <= X"40000278";
    when 16#114B# => romdata <= X"9607BFD0";
    when 16#114C# => romdata <= X"80A23FFF";
    when 16#114D# => romdata <= X"228001F4";
    when 16#114E# => romdata <= X"C416600C";
    when 16#114F# => romdata <= X"82020010";
    when 16#1150# => romdata <= X"80A0401D";
    when 16#1151# => romdata <= X"148001BA";
    when 16#1152# => romdata <= X"80A74001";
    when 16#1153# => romdata <= X"12BFFFF0";
    when 16#1154# => romdata <= X"AC05A004";
    when 16#1155# => romdata <= X"A0100015";
    when 16#1156# => romdata <= X"AA10001B";
    when 16#1157# => romdata <= X"F607B910";
    when 16#1158# => romdata <= X"80A76000";
    when 16#1159# => romdata <= X"12800192";
    when 16#115A# => romdata <= X"AC102000";
    when 16#115B# => romdata <= X"C027B910";
    when 16#115C# => romdata <= X"10BFFC80";
    when 16#115D# => romdata <= X"C027B908";
    when 16#115E# => romdata <= X"EE240000";
    when 16#115F# => romdata <= X"A0042008";
    when 16#1160# => romdata <= X"C407BFB4";
    when 16#1161# => romdata <= X"82008001";
    when 16#1162# => romdata <= X"C227BFB4";
    when 16#1163# => romdata <= X"C207BFB0";
    when 16#1164# => romdata <= X"82006001";
    when 16#1165# => romdata <= X"80A06007";
    when 16#1166# => romdata <= X"148000A6";
    when 16#1167# => romdata <= X"C227BFB0";
    when 16#1168# => romdata <= X"82102001";
    when 16#1169# => romdata <= X"EA07BFF4";
    when 16#116A# => romdata <= X"C2242004";
    when 16#116B# => romdata <= X"03100032";
    when 16#116C# => romdata <= X"82106050";
    when 16#116D# => romdata <= X"C407BFB4";
    when 16#116E# => romdata <= X"C2240000";
    when 16#116F# => romdata <= X"C207BFB0";
    when 16#1170# => romdata <= X"82006001";
    when 16#1171# => romdata <= X"8400A001";
    when 16#1172# => romdata <= X"C227BFB0";
    when 16#1173# => romdata <= X"C427BFB4";
    when 16#1174# => romdata <= X"80A06007";
    when 16#1175# => romdata <= X"1480008F";
    when 16#1176# => romdata <= X"A0042008";
    when 16#1177# => romdata <= X"C207BFF4";
    when 16#1178# => romdata <= X"C607B8F4";
    when 16#1179# => romdata <= X"8420C001";
    when 16#117A# => romdata <= X"C4242004";
    when 16#117B# => romdata <= X"AA05C015";
    when 16#117C# => romdata <= X"EA240000";
    when 16#117D# => romdata <= X"C407BFB4";
    when 16#117E# => romdata <= X"84208001";
    when 16#117F# => romdata <= X"C207BFB0";
    when 16#1180# => romdata <= X"10BFFDDB";
    when 16#1181# => romdata <= X"82006001";
    when 16#1182# => romdata <= X"EA242004";
    when 16#1183# => romdata <= X"C407B90C";
    when 16#1184# => romdata <= X"C4240000";
    when 16#1185# => romdata <= X"C207BFB4";
    when 16#1186# => romdata <= X"AA004015";
    when 16#1187# => romdata <= X"C207BFB0";
    when 16#1188# => romdata <= X"82006001";
    when 16#1189# => romdata <= X"EA27BFB4";
    when 16#118A# => romdata <= X"C227BFB0";
    when 16#118B# => romdata <= X"80A06007";
    when 16#118C# => romdata <= X"04800008";
    when 16#118D# => romdata <= X"A0042008";
    when 16#118E# => romdata <= X"90100019";
    when 16#118F# => romdata <= X"7FFFFAC5";
    when 16#1190# => romdata <= X"9207BFAC";
    when 16#1191# => romdata <= X"80A22000";
    when 16#1192# => romdata <= X"12BFFD3F";
    when 16#1193# => romdata <= X"A0100013";
    when 16#1194# => romdata <= X"808D2001";
    when 16#1195# => romdata <= X"02BFFB9B";
    when 16#1196# => romdata <= X"808D2004";
    when 16#1197# => romdata <= X"82102001";
    when 16#1198# => romdata <= X"C2242004";
    when 16#1199# => romdata <= X"03100032";
    when 16#119A# => romdata <= X"82106050";
    when 16#119B# => romdata <= X"C407BFB4";
    when 16#119C# => romdata <= X"C2240000";
    when 16#119D# => romdata <= X"C207BFB0";
    when 16#119E# => romdata <= X"82006001";
    when 16#119F# => romdata <= X"10BFFDBD";
    when 16#11A0# => romdata <= X"8400A001";
    when 16#11A1# => romdata <= X"80A5A000";
    when 16#11A2# => romdata <= X"22BFFEFB";
    when 16#11A3# => romdata <= X"AC102001";
    when 16#11A4# => romdata <= X"10BFFEFA";
    when 16#11A5# => romdata <= X"808D2008";
    when 16#11A6# => romdata <= X"90100019";
    when 16#11A7# => romdata <= X"7FFFFAAD";
    when 16#11A8# => romdata <= X"9207BFAC";
    when 16#11A9# => romdata <= X"80A22000";
    when 16#11AA# => romdata <= X"12BFFD27";
    when 16#11AB# => romdata <= X"A0100013";
    when 16#11AC# => romdata <= X"10BFFCEA";
    when 16#11AD# => romdata <= X"C207BFF4";
    when 16#11AE# => romdata <= X"84102004";
    when 16#11AF# => romdata <= X"2F100032";
    when 16#11B0# => romdata <= X"C22FBFFF";
    when 16#11B1# => romdata <= X"C427B910";
    when 16#11B2# => romdata <= X"BA102003";
    when 16#11B3# => romdata <= X"AE15E020";
    when 16#11B4# => romdata <= X"C027B908";
    when 16#11B5# => romdata <= X"10BFFC2E";
    when 16#11B6# => romdata <= X"AC102000";
    when 16#11B7# => romdata <= X"82102001";
    when 16#11B8# => romdata <= X"C2242004";
    when 16#11B9# => romdata <= X"03100032";
    when 16#11BA# => romdata <= X"82106048";
    when 16#11BB# => romdata <= X"C407BFB4";
    when 16#11BC# => romdata <= X"C2240000";
    when 16#11BD# => romdata <= X"C207BFB0";
    when 16#11BE# => romdata <= X"82006001";
    when 16#11BF# => romdata <= X"8400A001";
    when 16#11C0# => romdata <= X"C227BFB0";
    when 16#11C1# => romdata <= X"C427BFB4";
    when 16#11C2# => romdata <= X"80A06007";
    when 16#11C3# => romdata <= X"14800051";
    when 16#11C4# => romdata <= X"A0042008";
    when 16#11C5# => romdata <= X"C207BFF4";
    when 16#11C6# => romdata <= X"80A06000";
    when 16#11C7# => romdata <= X"02800030";
    when 16#11C8# => romdata <= X"C607B8F4";
    when 16#11C9# => romdata <= X"82102001";
    when 16#11CA# => romdata <= X"C2242004";
    when 16#11CB# => romdata <= X"C207B8E8";
    when 16#11CC# => romdata <= X"C2240000";
    when 16#11CD# => romdata <= X"C407BFB0";
    when 16#11CE# => romdata <= X"C607BFB4";
    when 16#11CF# => romdata <= X"8400A001";
    when 16#11D0# => romdata <= X"8600E001";
    when 16#11D1# => romdata <= X"C427BFB0";
    when 16#11D2# => romdata <= X"C627BFB4";
    when 16#11D3# => romdata <= X"80A0A007";
    when 16#11D4# => romdata <= X"14800164";
    when 16#11D5# => romdata <= X"82042008";
    when 16#11D6# => romdata <= X"EA07BFF4";
    when 16#11D7# => romdata <= X"AA200015";
    when 16#11D8# => romdata <= X"80A56000";
    when 16#11D9# => romdata <= X"048000F5";
    when 16#11DA# => romdata <= X"80A56010";
    when 16#11DB# => romdata <= X"048000E1";
    when 16#11DC# => romdata <= X"E227B90C";
    when 16#11DD# => romdata <= X"BA102010";
    when 16#11DE# => romdata <= X"10800006";
    when 16#11DF# => romdata <= X"A007BFAC";
    when 16#11E0# => romdata <= X"AA057FF0";
    when 16#11E1# => romdata <= X"80A56010";
    when 16#11E2# => romdata <= X"248000DB";
    when 16#11E3# => romdata <= X"EA206004";
    when 16#11E4# => romdata <= X"FA206004";
    when 16#11E5# => romdata <= X"E2204000";
    when 16#11E6# => romdata <= X"82006008";
    when 16#11E7# => romdata <= X"C407BFB0";
    when 16#11E8# => romdata <= X"C607BFB4";
    when 16#11E9# => romdata <= X"8400A001";
    when 16#11EA# => romdata <= X"8600E010";
    when 16#11EB# => romdata <= X"C427BFB0";
    when 16#11EC# => romdata <= X"80A0A007";
    when 16#11ED# => romdata <= X"04BFFFF3";
    when 16#11EE# => romdata <= X"C627BFB4";
    when 16#11EF# => romdata <= X"90100019";
    when 16#11F0# => romdata <= X"7FFFFA64";
    when 16#11F1# => romdata <= X"92100010";
    when 16#11F2# => romdata <= X"80A22000";
    when 16#11F3# => romdata <= X"12BFFCDE";
    when 16#11F4# => romdata <= X"82100013";
    when 16#11F5# => romdata <= X"10BFFFEC";
    when 16#11F6# => romdata <= X"AA057FF0";
    when 16#11F7# => romdata <= X"80A0E000";
    when 16#11F8# => romdata <= X"02BFFB38";
    when 16#11F9# => romdata <= X"808D2004";
    when 16#11FA# => romdata <= X"10BFFFD0";
    when 16#11FB# => romdata <= X"82102001";
    when 16#11FC# => romdata <= X"90100019";
    when 16#11FD# => romdata <= X"7FFFFA57";
    when 16#11FE# => romdata <= X"9207BFAC";
    when 16#11FF# => romdata <= X"80A22000";
    when 16#1200# => romdata <= X"12BFFCD1";
    when 16#1201# => romdata <= X"A0100013";
    when 16#1202# => romdata <= X"10BFFD8E";
    when 16#1203# => romdata <= X"EA07BFF4";
    when 16#1204# => romdata <= X"90100019";
    when 16#1205# => romdata <= X"7FFFFA4F";
    when 16#1206# => romdata <= X"9207BFAC";
    when 16#1207# => romdata <= X"80A22000";
    when 16#1208# => romdata <= X"12BFFCC9";
    when 16#1209# => romdata <= X"A0100013";
    when 16#120A# => romdata <= X"10BFFF6E";
    when 16#120B# => romdata <= X"C207BFF4";
    when 16#120C# => romdata <= X"90100019";
    when 16#120D# => romdata <= X"7FFFFA47";
    when 16#120E# => romdata <= X"9207BFAC";
    when 16#120F# => romdata <= X"80A22000";
    when 16#1210# => romdata <= X"12BFFCC1";
    when 16#1211# => romdata <= X"A0100013";
    when 16#1212# => romdata <= X"10BFFF57";
    when 16#1213# => romdata <= X"82102001";
    when 16#1214# => romdata <= X"90100019";
    when 16#1215# => romdata <= X"7FFFFA3F";
    when 16#1216# => romdata <= X"9207BFAC";
    when 16#1217# => romdata <= X"80A22000";
    when 16#1218# => romdata <= X"12BFFCB9";
    when 16#1219# => romdata <= X"A0100013";
    when 16#121A# => romdata <= X"10BFFFAC";
    when 16#121B# => romdata <= X"C207BFF4";
    when 16#121C# => romdata <= X"C027B908";
    when 16#121D# => romdata <= X"4000136A";
    when 16#121E# => romdata <= X"AC102000";
    when 16#121F# => romdata <= X"82380008";
    when 16#1220# => romdata <= X"BA100008";
    when 16#1221# => romdata <= X"8338601F";
    when 16#1222# => romdata <= X"820A0001";
    when 16#1223# => romdata <= X"10BFFBB9";
    when 16#1224# => romdata <= X"C227B910";
    when 16#1225# => romdata <= X"C207BFB4";
    when 16#1226# => romdata <= X"80A06000";
    when 16#1227# => romdata <= X"12800005";
    when 16#1228# => romdata <= X"90100019";
    when 16#1229# => romdata <= X"C027BFB0";
    when 16#122A# => romdata <= X"10BFFCAE";
    when 16#122B# => romdata <= X"C216600C";
    when 16#122C# => romdata <= X"7FFFFA28";
    when 16#122D# => romdata <= X"9207BFAC";
    when 16#122E# => romdata <= X"80A22000";
    when 16#122F# => romdata <= X"32BFFCA9";
    when 16#1230# => romdata <= X"C216600C";
    when 16#1231# => romdata <= X"C027BFB0";
    when 16#1232# => romdata <= X"10BFFCA6";
    when 16#1233# => romdata <= X"C216600C";
    when 16#1234# => romdata <= X"10BFFE69";
    when 16#1235# => romdata <= X"AC102006";
    when 16#1236# => romdata <= X"EA0E8000";
    when 16#1237# => romdata <= X"A8152010";
    when 16#1238# => romdata <= X"10BFFA81";
    when 16#1239# => romdata <= X"AB2D6018";
    when 16#123A# => romdata <= X"400012FC";
    when 16#123B# => romdata <= X"D01FB8F8";
    when 16#123C# => romdata <= X"80A22000";
    when 16#123D# => romdata <= X"128000A7";
    when 16#123E# => romdata <= X"86102003";
    when 16#123F# => romdata <= X"A8152100";
    when 16#1240# => romdata <= X"80A56066";
    when 16#1241# => romdata <= X"BA100016";
    when 16#1242# => romdata <= X"02800007";
    when 16#1243# => romdata <= X"96102003";
    when 16#1244# => romdata <= X"80A56045";
    when 16#1245# => romdata <= X"02800100";
    when 16#1246# => romdata <= X"80A56065";
    when 16#1247# => romdata <= X"028000FE";
    when 16#1248# => romdata <= X"96102002";
    when 16#1249# => romdata <= X"D11FB8F8";
    when 16#124A# => romdata <= X"D13FBFB8";
    when 16#124B# => romdata <= X"C02FB90C";
    when 16#124C# => romdata <= X"C207BFB8";
    when 16#124D# => romdata <= X"80A06000";
    when 16#124E# => romdata <= X"0680011D";
    when 16#124F# => romdata <= X"95A00028";
    when 16#1250# => romdata <= X"8207BFEC";
    when 16#1251# => romdata <= X"D007A044";
    when 16#1252# => romdata <= X"C223A05C";
    when 16#1253# => romdata <= X"D207B910";
    when 16#1254# => romdata <= X"8207BFE8";
    when 16#1255# => romdata <= X"D407B914";
    when 16#1256# => romdata <= X"C223A060";
    when 16#1257# => romdata <= X"9810001D";
    when 16#1258# => romdata <= X"400003B8";
    when 16#1259# => romdata <= X"9A07BFF4";
    when 16#125A# => romdata <= X"80A56047";
    when 16#125B# => romdata <= X"028000C2";
    when 16#125C# => romdata <= X"AE100008";
    when 16#125D# => romdata <= X"80A56067";
    when 16#125E# => romdata <= X"028000C0";
    when 16#125F# => romdata <= X"808D2001";
    when 16#1260# => romdata <= X"03100032";
    when 16#1261# => romdata <= X"80A56066";
    when 16#1262# => romdata <= X"8405C01D";
    when 16#1263# => romdata <= X"0280010E";
    when 16#1264# => romdata <= X"82106060";
    when 16#1265# => romdata <= X"D1184000";
    when 16#1266# => romdata <= X"D51FB910";
    when 16#1267# => romdata <= X"81AA8A48";
    when 16#1268# => romdata <= X"01000000";
    when 16#1269# => romdata <= X"038000B9";
    when 16#126A# => romdata <= X"C807BFE8";
    when 16#126B# => romdata <= X"C427BFE8";
    when 16#126C# => romdata <= X"821D6067";
    when 16#126D# => romdata <= X"84208017";
    when 16#126E# => romdata <= X"80A00001";
    when 16#126F# => romdata <= X"82603FFF";
    when 16#1270# => romdata <= X"80A56047";
    when 16#1271# => romdata <= X"02800005";
    when 16#1272# => romdata <= X"C427B8F4";
    when 16#1273# => romdata <= X"80A06000";
    when 16#1274# => romdata <= X"0280009C";
    when 16#1275# => romdata <= X"80A56065";
    when 16#1276# => romdata <= X"FA07BFF4";
    when 16#1277# => romdata <= X"80A77FFD";
    when 16#1278# => romdata <= X"06800006";
    when 16#1279# => romdata <= X"80A06000";
    when 16#127A# => romdata <= X"80A5801D";
    when 16#127B# => romdata <= X"1680009A";
    when 16#127C# => romdata <= X"C607B8F4";
    when 16#127D# => romdata <= X"80A06000";
    when 16#127E# => romdata <= X"AA102045";
    when 16#127F# => romdata <= X"02800004";
    when 16#1280# => romdata <= X"82102045";
    when 16#1281# => romdata <= X"82102065";
    when 16#1282# => romdata <= X"AA102065";
    when 16#1283# => romdata <= X"BA077FFF";
    when 16#1284# => romdata <= X"C22FBFE0";
    when 16#1285# => romdata <= X"80A76000";
    when 16#1286# => romdata <= X"06800108";
    when 16#1287# => romdata <= X"FA27BFF4";
    when 16#1288# => romdata <= X"8210202B";
    when 16#1289# => romdata <= X"C22FBFE1";
    when 16#128A# => romdata <= X"80A76009";
    when 16#128B# => romdata <= X"148000BD";
    when 16#128C# => romdata <= X"8207BFA8";
    when 16#128D# => romdata <= X"BA076030";
    when 16#128E# => romdata <= X"82102030";
    when 16#128F# => romdata <= X"C22FBFE2";
    when 16#1290# => romdata <= X"FA2FBFE3";
    when 16#1291# => romdata <= X"8407BFE4";
    when 16#1292# => romdata <= X"C207B8F4";
    when 16#1293# => romdata <= X"80A06001";
    when 16#1294# => romdata <= X"8207BFE0";
    when 16#1295# => romdata <= X"82208001";
    when 16#1296# => romdata <= X"C407B8F4";
    when 16#1297# => romdata <= X"C227B8F0";
    when 16#1298# => romdata <= X"04800011";
    when 16#1299# => romdata <= X"BA004002";
    when 16#129A# => romdata <= X"BA076001";
    when 16#129B# => romdata <= X"C40FB90C";
    when 16#129C# => romdata <= X"8088A0FF";
    when 16#129D# => romdata <= X"02800019";
    when 16#129E# => romdata <= X"8238001D";
    when 16#129F# => romdata <= X"8210202D";
    when 16#12A0# => romdata <= X"C027B908";
    when 16#12A1# => romdata <= X"C22FBFFF";
    when 16#12A2# => romdata <= X"AC102000";
    when 16#12A3# => romdata <= X"8238001D";
    when 16#12A4# => romdata <= X"8338601F";
    when 16#12A5# => romdata <= X"820F4001";
    when 16#12A6# => romdata <= X"82006001";
    when 16#12A7# => romdata <= X"10BFFB3C";
    when 16#12A8# => romdata <= X"C227B910";
    when 16#12A9# => romdata <= X"808D2001";
    when 16#12AA# => romdata <= X"02BFFFF2";
    when 16#12AB# => romdata <= X"C40FB90C";
    when 16#12AC# => romdata <= X"10BFFFF0";
    when 16#12AD# => romdata <= X"BA076001";
    when 16#12AE# => romdata <= X"90100019";
    when 16#12AF# => romdata <= X"7FFFF9A5";
    when 16#12B0# => romdata <= X"9207BFAC";
    when 16#12B1# => romdata <= X"80A22000";
    when 16#12B2# => romdata <= X"12BFFC1F";
    when 16#12B3# => romdata <= X"A0100013";
    when 16#12B4# => romdata <= X"10BFFBF7";
    when 16#12B5# => romdata <= X"C207B8F4";
    when 16#12B6# => romdata <= X"C027B908";
    when 16#12B7# => romdata <= X"8338601F";
    when 16#12B8# => romdata <= X"AC102000";
    when 16#12B9# => romdata <= X"820F4001";
    when 16#12BA# => romdata <= X"10BFFB22";
    when 16#12BB# => romdata <= X"C227B910";
    when 16#12BC# => romdata <= X"EA206004";
    when 16#12BD# => romdata <= X"C407B90C";
    when 16#12BE# => romdata <= X"C4204000";
    when 16#12BF# => romdata <= X"C407BFB4";
    when 16#12C0# => romdata <= X"AA008015";
    when 16#12C1# => romdata <= X"C407BFB0";
    when 16#12C2# => romdata <= X"8400A001";
    when 16#12C3# => romdata <= X"EA27BFB4";
    when 16#12C4# => romdata <= X"C427BFB0";
    when 16#12C5# => romdata <= X"80A0A007";
    when 16#12C6# => romdata <= X"04800008";
    when 16#12C7# => romdata <= X"82006008";
    when 16#12C8# => romdata <= X"90100019";
    when 16#12C9# => romdata <= X"7FFFF98B";
    when 16#12CA# => romdata <= X"9207BFAC";
    when 16#12CB# => romdata <= X"80A22000";
    when 16#12CC# => romdata <= X"12BFFC05";
    when 16#12CD# => romdata <= X"82100013";
    when 16#12CE# => romdata <= X"C607B8F4";
    when 16#12CF# => romdata <= X"C6206004";
    when 16#12D0# => romdata <= X"EE204000";
    when 16#12D1# => romdata <= X"A0006008";
    when 16#12D2# => romdata <= X"C407BFB4";
    when 16#12D3# => romdata <= X"C207BFB0";
    when 16#12D4# => romdata <= X"82006001";
    when 16#12D5# => romdata <= X"84008003";
    when 16#12D6# => romdata <= X"C227BFB0";
    when 16#12D7# => romdata <= X"80A06007";
    when 16#12D8# => romdata <= X"04BFFA57";
    when 16#12D9# => romdata <= X"C427BFB4";
    when 16#12DA# => romdata <= X"10BFFC88";
    when 16#12DB# => romdata <= X"90100019";
    when 16#12DC# => romdata <= X"82102006";
    when 16#12DD# => romdata <= X"2F100032";
    when 16#12DE# => romdata <= X"C227B910";
    when 16#12DF# => romdata <= X"BA102006";
    when 16#12E0# => romdata <= X"AE15E058";
    when 16#12E1# => romdata <= X"C027B908";
    when 16#12E2# => romdata <= X"10BFF9E7";
    when 16#12E3# => romdata <= X"AC102000";
    when 16#12E4# => romdata <= X"2F100032";
    when 16#12E5# => romdata <= X"C627B910";
    when 16#12E6# => romdata <= X"BA102003";
    when 16#12E7# => romdata <= X"C027B908";
    when 16#12E8# => romdata <= X"AE15E040";
    when 16#12E9# => romdata <= X"10BFFAF3";
    when 16#12EA# => romdata <= X"AC102000";
    when 16#12EB# => romdata <= X"D007A044";
    when 16#12EC# => romdata <= X"7FFFF73D";
    when 16#12ED# => romdata <= X"92076001";
    when 16#12EE# => romdata <= X"AC922000";
    when 16#12EF# => romdata <= X"02800051";
    when 16#12F0# => romdata <= X"94102008";
    when 16#12F1# => romdata <= X"92102000";
    when 16#12F2# => romdata <= X"40000CB8";
    when 16#12F3# => romdata <= X"9007BFD0";
    when 16#12F4# => romdata <= X"D007A044";
    when 16#12F5# => romdata <= X"92100016";
    when 16#12F6# => romdata <= X"9807BFD0";
    when 16#12F7# => romdata <= X"9407BFF0";
    when 16#12F8# => romdata <= X"400000ED";
    when 16#12F9# => romdata <= X"9610001D";
    when 16#12FA# => romdata <= X"80A74008";
    when 16#12FB# => romdata <= X"128000B8";
    when 16#12FC# => romdata <= X"8238001D";
    when 16#12FD# => romdata <= X"C02D801D";
    when 16#12FE# => romdata <= X"AE100016";
    when 16#12FF# => romdata <= X"8338601F";
    when 16#1300# => romdata <= X"C027B908";
    when 16#1301# => romdata <= X"820F4001";
    when 16#1302# => romdata <= X"10BFFADA";
    when 16#1303# => romdata <= X"C227B910";
    when 16#1304# => romdata <= X"80886200";
    when 16#1305# => romdata <= X"12BFFBDD";
    when 16#1306# => romdata <= X"90066058";
    when 16#1307# => romdata <= X"400017B3";
    when 16#1308# => romdata <= X"B0103FFF";
    when 16#1309# => romdata <= X"81C7E008";
    when 16#130A# => romdata <= X"81E80000";
    when 16#130B# => romdata <= X"BA100010";
    when 16#130C# => romdata <= X"A0100015";
    when 16#130D# => romdata <= X"AA10001B";
    when 16#130E# => romdata <= X"10BFFE4A";
    when 16#130F# => romdata <= X"F607B910";
    when 16#1310# => romdata <= X"04800058";
    when 16#1311# => romdata <= X"80A56066";
    when 16#1312# => romdata <= X"0280008B";
    when 16#1313# => romdata <= X"FA07BFF4";
    when 16#1314# => romdata <= X"C607B8F4";
    when 16#1315# => romdata <= X"80A0C01D";
    when 16#1316# => romdata <= X"14800063";
    when 16#1317# => romdata <= X"80A76000";
    when 16#1318# => romdata <= X"808D2001";
    when 16#1319# => romdata <= X"02BFFF82";
    when 16#131A# => romdata <= X"AA102067";
    when 16#131B# => romdata <= X"10BFFF80";
    when 16#131C# => romdata <= X"BA076001";
    when 16#131D# => romdata <= X"808D2001";
    when 16#131E# => romdata <= X"12BFFF43";
    when 16#131F# => romdata <= X"03100032";
    when 16#1320# => romdata <= X"10BFFF4C";
    when 16#1321# => romdata <= X"C407BFE8";
    when 16#1322# => romdata <= X"80A08004";
    when 16#1323# => romdata <= X"82100004";
    when 16#1324# => romdata <= X"0880008D";
    when 16#1325# => romdata <= X"86102030";
    when 16#1326# => romdata <= X"C6284000";
    when 16#1327# => romdata <= X"82006001";
    when 16#1328# => romdata <= X"80A08001";
    when 16#1329# => romdata <= X"18BFFFFD";
    when 16#132A# => romdata <= X"C227BFE8";
    when 16#132B# => romdata <= X"10BFFF42";
    when 16#132C# => romdata <= X"821D6067";
    when 16#132D# => romdata <= X"D007A044";
    when 16#132E# => romdata <= X"92102000";
    when 16#132F# => romdata <= X"9407BFF0";
    when 16#1330# => romdata <= X"96102000";
    when 16#1331# => romdata <= X"400000B4";
    when 16#1332# => romdata <= X"9807BFD0";
    when 16#1333# => romdata <= X"80A23FFF";
    when 16#1334# => romdata <= X"0280000C";
    when 16#1335# => romdata <= X"BA100008";
    when 16#1336# => romdata <= X"10BFFE22";
    when 16#1337# => romdata <= X"EE27BFF0";
    when 16#1338# => romdata <= X"90100019";
    when 16#1339# => romdata <= X"7FFFF91B";
    when 16#133A# => romdata <= X"9207BFAC";
    when 16#133B# => romdata <= X"80A22000";
    when 16#133C# => romdata <= X"12BFFB95";
    when 16#133D# => romdata <= X"82100013";
    when 16#133E# => romdata <= X"10BFFE99";
    when 16#133F# => romdata <= X"EA07BFF4";
    when 16#1340# => romdata <= X"C416600C";
    when 16#1341# => romdata <= X"8410A040";
    when 16#1342# => romdata <= X"82100002";
    when 16#1343# => romdata <= X"10BFFB95";
    when 16#1344# => romdata <= X"C436600C";
    when 16#1345# => romdata <= X"BA05A001";
    when 16#1346# => romdata <= X"10BFFF03";
    when 16#1347# => romdata <= X"96102002";
    when 16#1348# => romdata <= X"AC100001";
    when 16#1349# => romdata <= X"C227B8E4";
    when 16#134A# => romdata <= X"9010001D";
    when 16#134B# => romdata <= X"9210200A";
    when 16#134C# => romdata <= X"4000142A";
    when 16#134D# => romdata <= X"AC05BFFF";
    when 16#134E# => romdata <= X"84022030";
    when 16#134F# => romdata <= X"9210200A";
    when 16#1350# => romdata <= X"9010001D";
    when 16#1351# => romdata <= X"40001379";
    when 16#1352# => romdata <= X"C42D8000";
    when 16#1353# => romdata <= X"C207B8E4";
    when 16#1354# => romdata <= X"80A22009";
    when 16#1355# => romdata <= X"14BFFFF4";
    when 16#1356# => romdata <= X"BA100008";
    when 16#1357# => romdata <= X"88022030";
    when 16#1358# => romdata <= X"8405BFFF";
    when 16#1359# => romdata <= X"86100016";
    when 16#135A# => romdata <= X"C82DBFFF";
    when 16#135B# => romdata <= X"80A04002";
    when 16#135C# => romdata <= X"18800006";
    when 16#135D# => romdata <= X"8407BFE2";
    when 16#135E# => romdata <= X"10BFFF35";
    when 16#135F# => romdata <= X"C207B8F4";
    when 16#1360# => romdata <= X"C808C000";
    when 16#1361# => romdata <= X"8600E001";
    when 16#1362# => romdata <= X"C8288000";
    when 16#1363# => romdata <= X"80A04003";
    when 16#1364# => romdata <= X"18BFFFFC";
    when 16#1365# => romdata <= X"8400A001";
    when 16#1366# => romdata <= X"10BFFF2D";
    when 16#1367# => romdata <= X"C207B8F4";
    when 16#1368# => romdata <= X"FA07BFF4";
    when 16#1369# => romdata <= X"10BFFF1A";
    when 16#136A# => romdata <= X"82100015";
    when 16#136B# => romdata <= X"97A00029";
    when 16#136C# => romdata <= X"95A000AA";
    when 16#136D# => romdata <= X"8210202D";
    when 16#136E# => romdata <= X"D53FB910";
    when 16#136F# => romdata <= X"10BFFEE1";
    when 16#1370# => romdata <= X"C22FB90C";
    when 16#1371# => romdata <= X"C24DC000";
    when 16#1372# => romdata <= X"80A06030";
    when 16#1373# => romdata <= X"0280000E";
    when 16#1374# => romdata <= X"03100032";
    when 16#1375# => romdata <= X"FA07BFF4";
    when 16#1376# => romdata <= X"8400801D";
    when 16#1377# => romdata <= X"10BFFEEE";
    when 16#1378# => romdata <= X"82106060";
    when 16#1379# => romdata <= X"82102002";
    when 16#137A# => romdata <= X"04800003";
    when 16#137B# => romdata <= X"BA20401D";
    when 16#137C# => romdata <= X"BA102001";
    when 16#137D# => romdata <= X"C207B8F4";
    when 16#137E# => romdata <= X"BA074001";
    when 16#137F# => romdata <= X"10BFFF1C";
    when 16#1380# => romdata <= X"AA102067";
    when 16#1381# => romdata <= X"07100032";
    when 16#1382# => romdata <= X"D51FB910";
    when 16#1383# => romdata <= X"8610E060";
    when 16#1384# => romdata <= X"D118C000";
    when 16#1385# => romdata <= X"81AA8A48";
    when 16#1386# => romdata <= X"01000000";
    when 16#1387# => romdata <= X"1380000B";
    when 16#1388# => romdata <= X"82100003";
    when 16#1389# => romdata <= X"86102001";
    when 16#138A# => romdata <= X"BA20C01D";
    when 16#138B# => romdata <= X"FA27BFF4";
    when 16#138C# => romdata <= X"10BFFED9";
    when 16#138D# => romdata <= X"8400801D";
    when 16#138E# => romdata <= X"8210202D";
    when 16#138F# => romdata <= X"BA20001D";
    when 16#1390# => romdata <= X"10BFFEFA";
    when 16#1391# => romdata <= X"C22FBFE1";
    when 16#1392# => romdata <= X"FA07BFF4";
    when 16#1393# => romdata <= X"10BFFED2";
    when 16#1394# => romdata <= X"8400801D";
    when 16#1395# => romdata <= X"EC06C000";
    when 16#1396# => romdata <= X"80A5A000";
    when 16#1397# => romdata <= X"16BFFC70";
    when 16#1398# => romdata <= X"B606E004";
    when 16#1399# => romdata <= X"EA0E8000";
    when 16#139A# => romdata <= X"AB2D6018";
    when 16#139B# => romdata <= X"10BFF91E";
    when 16#139C# => romdata <= X"AC103FFF";
    when 16#139D# => romdata <= X"80A76000";
    when 16#139E# => romdata <= X"0480000B";
    when 16#139F# => romdata <= X"80A5A000";
    when 16#13A0# => romdata <= X"32800006";
    when 16#13A1# => romdata <= X"BA076001";
    when 16#13A2# => romdata <= X"808D2001";
    when 16#13A3# => romdata <= X"02BFFEF9";
    when 16#13A4# => romdata <= X"C40FB90C";
    when 16#13A5# => romdata <= X"BA076001";
    when 16#13A6# => romdata <= X"AA102066";
    when 16#13A7# => romdata <= X"10BFFEF4";
    when 16#13A8# => romdata <= X"BA074016";
    when 16#13A9# => romdata <= X"12800006";
    when 16#13AA# => romdata <= X"BA05A002";
    when 16#13AB# => romdata <= X"808D2001";
    when 16#13AC# => romdata <= X"02BFFEEF";
    when 16#13AD# => romdata <= X"BA102001";
    when 16#13AE# => romdata <= X"BA05A002";
    when 16#13AF# => romdata <= X"10BFFEEC";
    when 16#13B0# => romdata <= X"AA102066";
    when 16#13B1# => romdata <= X"10BFFEBB";
    when 16#13B2# => romdata <= X"84100004";
    when 16#13B3# => romdata <= X"C216600C";
    when 16#13B4# => romdata <= X"82106040";
    when 16#13B5# => romdata <= X"10BFFB1F";
    when 16#13B6# => romdata <= X"C236600C";
    when 16#13B7# => romdata <= X"03100032";
    when 16#13B8# => romdata <= X"84100008";
    when 16#13B9# => romdata <= X"D00062C8";
    when 16#13BA# => romdata <= X"82100009";
    when 16#13BB# => romdata <= X"9610000A";
    when 16#13BC# => romdata <= X"92100002";
    when 16#13BD# => romdata <= X"94100001";
    when 16#13BE# => romdata <= X"8213C000";
    when 16#13BF# => romdata <= X"7FFFF8A3";
    when 16#13C0# => romdata <= X"9E104000";
    when 16#13C1# => romdata <= X"01000000";
    when 16#13C2# => romdata <= X"9DE3BF90";
    when 16#13C3# => romdata <= X"80A66000";
    when 16#13C4# => romdata <= X"0280000F";
    when 16#13C5# => romdata <= X"A0100018";
    when 16#13C6# => romdata <= X"92100019";
    when 16#13C7# => romdata <= X"9410001A";
    when 16#13C8# => romdata <= X"90100018";
    when 16#13C9# => romdata <= X"40000077";
    when 16#13CA# => romdata <= X"9610001B";
    when 16#13CB# => romdata <= X"80A23FFF";
    when 16#13CC# => romdata <= X"12800005";
    when 16#13CD# => romdata <= X"B0100008";
    when 16#13CE# => romdata <= X"C026C000";
    when 16#13CF# => romdata <= X"8210208A";
    when 16#13D0# => romdata <= X"C2240000";
    when 16#13D1# => romdata <= X"81C7E008";
    when 16#13D2# => romdata <= X"81E80000";
    when 16#13D3# => romdata <= X"90100018";
    when 16#13D4# => romdata <= X"9207BFF0";
    when 16#13D5# => romdata <= X"94102000";
    when 16#13D6# => romdata <= X"4000006A";
    when 16#13D7# => romdata <= X"9610001B";
    when 16#13D8# => romdata <= X"10BFFFF4";
    when 16#13D9# => romdata <= X"80A23FFF";
    when 16#13DA# => romdata <= X"03100032";
    when 16#13DB# => romdata <= X"84100008";
    when 16#13DC# => romdata <= X"D00062C8";
    when 16#13DD# => romdata <= X"82100009";
    when 16#13DE# => romdata <= X"9610000A";
    when 16#13DF# => romdata <= X"92100002";
    when 16#13E0# => romdata <= X"94100001";
    when 16#13E1# => romdata <= X"8213C000";
    when 16#13E2# => romdata <= X"7FFFFFE0";
    when 16#13E3# => romdata <= X"9E104000";
    when 16#13E4# => romdata <= X"01000000";
    when 16#13E5# => romdata <= X"9DE3BF90";
    when 16#13E6# => romdata <= X"80A66000";
    when 16#13E7# => romdata <= X"02800049";
    when 16#13E8# => romdata <= X"A0100018";
    when 16#13E9# => romdata <= X"80A6E000";
    when 16#13EA# => romdata <= X"0280003D";
    when 16#13EB# => romdata <= X"E6068000";
    when 16#13EC# => romdata <= X"D404C000";
    when 16#13ED# => romdata <= X"A207BFF0";
    when 16#13EE# => romdata <= X"E8070000";
    when 16#13EF# => romdata <= X"EA072004";
    when 16#13F0# => romdata <= X"90100010";
    when 16#13F1# => romdata <= X"92100011";
    when 16#13F2# => romdata <= X"9610001C";
    when 16#13F3# => romdata <= X"7FFFFFCF";
    when 16#13F4# => romdata <= X"A4100019";
    when 16#13F5# => romdata <= X"80A23FFF";
    when 16#13F6# => romdata <= X"02800029";
    when 16#13F7# => romdata <= X"B0102000";
    when 16#13F8# => romdata <= X"8226C008";
    when 16#13F9# => romdata <= X"80A04018";
    when 16#13FA# => romdata <= X"2A80002A";
    when 16#13FB# => romdata <= X"EA272004";
    when 16#13FC# => romdata <= X"80A2001B";
    when 16#13FD# => romdata <= X"3A800027";
    when 16#13FE# => romdata <= X"EA272004";
    when 16#13FF# => romdata <= X"80A66000";
    when 16#1400# => romdata <= X"0280000F";
    when 16#1401# => romdata <= X"B0060008";
    when 16#1402# => romdata <= X"80A22000";
    when 16#1403# => romdata <= X"04800009";
    when 16#1404# => romdata <= X"82102000";
    when 16#1405# => romdata <= X"C40C4001";
    when 16#1406# => romdata <= X"C42C8001";
    when 16#1407# => romdata <= X"82006001";
    when 16#1408# => romdata <= X"80A20001";
    when 16#1409# => romdata <= X"32BFFFFD";
    when 16#140A# => romdata <= X"C40C4001";
    when 16#140B# => romdata <= X"A4048008";
    when 16#140C# => romdata <= X"C2068000";
    when 16#140D# => romdata <= X"82006004";
    when 16#140E# => romdata <= X"C2268000";
    when 16#140F# => romdata <= X"C204C000";
    when 16#1410# => romdata <= X"80A06000";
    when 16#1411# => romdata <= X"02800019";
    when 16#1412# => romdata <= X"80A6001B";
    when 16#1413# => romdata <= X"1A800012";
    when 16#1414# => romdata <= X"A604E004";
    when 16#1415# => romdata <= X"D404C000";
    when 16#1416# => romdata <= X"E8070000";
    when 16#1417# => romdata <= X"EA072004";
    when 16#1418# => romdata <= X"90100010";
    when 16#1419# => romdata <= X"92100011";
    when 16#141A# => romdata <= X"7FFFFFA8";
    when 16#141B# => romdata <= X"9610001C";
    when 16#141C# => romdata <= X"80A23FFF";
    when 16#141D# => romdata <= X"12BFFFDC";
    when 16#141E# => romdata <= X"8226C008";
    when 16#141F# => romdata <= X"8210208A";
    when 16#1420# => romdata <= X"C2240000";
    when 16#1421# => romdata <= X"C0270000";
    when 16#1422# => romdata <= X"81C7E008";
    when 16#1423# => romdata <= X"91E83FFF";
    when 16#1424# => romdata <= X"E8270000";
    when 16#1425# => romdata <= X"81C7E008";
    when 16#1426# => romdata <= X"81E80000";
    when 16#1427# => romdata <= X"B0102000";
    when 16#1428# => romdata <= X"81C7E008";
    when 16#1429# => romdata <= X"81E80000";
    when 16#142A# => romdata <= X"80A66000";
    when 16#142B# => romdata <= X"32800002";
    when 16#142C# => romdata <= X"C0268000";
    when 16#142D# => romdata <= X"C0270000";
    when 16#142E# => romdata <= X"81C7E008";
    when 16#142F# => romdata <= X"91EE3FFF";
    when 16#1430# => romdata <= X"E6068000";
    when 16#1431# => romdata <= X"10BFFFBB";
    when 16#1432# => romdata <= X"B6103FFF";
    when 16#1433# => romdata <= X"03100032";
    when 16#1434# => romdata <= X"86100008";
    when 16#1435# => romdata <= X"84100009";
    when 16#1436# => romdata <= X"D00062C8";
    when 16#1437# => romdata <= X"8210000A";
    when 16#1438# => romdata <= X"9810000B";
    when 16#1439# => romdata <= X"92100003";
    when 16#143A# => romdata <= X"94100002";
    when 16#143B# => romdata <= X"96100001";
    when 16#143C# => romdata <= X"8213C000";
    when 16#143D# => romdata <= X"7FFFFFA8";
    when 16#143E# => romdata <= X"9E104000";
    when 16#143F# => romdata <= X"01000000";
    when 16#1440# => romdata <= X"9DE3BFA0";
    when 16#1441# => romdata <= X"21100035";
    when 16#1442# => romdata <= X"40001145";
    when 16#1443# => romdata <= X"90142120";
    when 16#1444# => romdata <= X"80A22001";
    when 16#1445# => romdata <= X"08800027";
    when 16#1446# => romdata <= X"90142120";
    when 16#1447# => romdata <= X"13100032";
    when 16#1448# => romdata <= X"7FFFF525";
    when 16#1449# => romdata <= X"92126088";
    when 16#144A# => romdata <= X"80A22000";
    when 16#144B# => romdata <= X"12800012";
    when 16#144C# => romdata <= X"80A66000";
    when 16#144D# => romdata <= X"02800022";
    when 16#144E# => romdata <= X"80A6A07F";
    when 16#144F# => romdata <= X"2480001B";
    when 16#1450# => romdata <= X"F42E4000";
    when 16#1451# => romdata <= X"8206BF80";
    when 16#1452# => romdata <= X"80A0677F";
    when 16#1453# => romdata <= X"1880001E";
    when 16#1454# => romdata <= X"820EA03F";
    when 16#1455# => romdata <= X"B40EA7C0";
    when 16#1456# => romdata <= X"82107F80";
    when 16#1457# => romdata <= X"B53EA006";
    when 16#1458# => romdata <= X"B416BFC0";
    when 16#1459# => romdata <= X"C22E6001";
    when 16#145A# => romdata <= X"F42E4000";
    when 16#145B# => romdata <= X"81C7E008";
    when 16#145C# => romdata <= X"91E82002";
    when 16#145D# => romdata <= X"90142120";
    when 16#145E# => romdata <= X"13100032";
    when 16#145F# => romdata <= X"7FFFF50E";
    when 16#1460# => romdata <= X"92126090";
    when 16#1461# => romdata <= X"80A22000";
    when 16#1462# => romdata <= X"12800058";
    when 16#1463# => romdata <= X"80A66000";
    when 16#1464# => romdata <= X"0280000B";
    when 16#1465# => romdata <= X"833EA008";
    when 16#1466# => romdata <= X"848860FF";
    when 16#1467# => romdata <= X"12800041";
    when 16#1468# => romdata <= X"86006020";
    when 16#1469# => romdata <= X"F42E4000";
    when 16#146A# => romdata <= X"81C7E008";
    when 16#146B# => romdata <= X"91E82001";
    when 16#146C# => romdata <= X"80A66000";
    when 16#146D# => romdata <= X"32BFFFFD";
    when 16#146E# => romdata <= X"F42E4000";
    when 16#146F# => romdata <= X"81C7E008";
    when 16#1470# => romdata <= X"91E82000";
    when 16#1471# => romdata <= X"8406B800";
    when 16#1472# => romdata <= X"0300003D";
    when 16#1473# => romdata <= X"821063FF";
    when 16#1474# => romdata <= X"80A08001";
    when 16#1475# => romdata <= X"08800074";
    when 16#1476# => romdata <= X"053FFFC0";
    when 16#1477# => romdata <= X"030007BF";
    when 16#1478# => romdata <= X"84068002";
    when 16#1479# => romdata <= X"821063FF";
    when 16#147A# => romdata <= X"80A08001";
    when 16#147B# => romdata <= X"18800012";
    when 16#147C# => romdata <= X"880EA03F";
    when 16#147D# => romdata <= X"8736A012";
    when 16#147E# => romdata <= X"88113F80";
    when 16#147F# => romdata <= X"8608E007";
    when 16#1480# => romdata <= X"8536A00C";
    when 16#1481# => romdata <= X"8610FFF0";
    when 16#1482# => romdata <= X"8408A03F";
    when 16#1483# => romdata <= X"820EAFC0";
    when 16#1484# => romdata <= X"8410BF80";
    when 16#1485# => romdata <= X"83386006";
    when 16#1486# => romdata <= X"82107F80";
    when 16#1487# => romdata <= X"C82E6003";
    when 16#1488# => romdata <= X"C62E4000";
    when 16#1489# => romdata <= X"C42E6001";
    when 16#148A# => romdata <= X"C22E6002";
    when 16#148B# => romdata <= X"81C7E008";
    when 16#148C# => romdata <= X"91E82004";
    when 16#148D# => romdata <= X"053FF800";
    when 16#148E# => romdata <= X"0300F7FF";
    when 16#148F# => romdata <= X"84068002";
    when 16#1490# => romdata <= X"821063FF";
    when 16#1491# => romdata <= X"80A08001";
    when 16#1492# => romdata <= X"1880006E";
    when 16#1493# => romdata <= X"9A0EA03F";
    when 16#1494# => romdata <= X"8936A018";
    when 16#1495# => romdata <= X"9A137F80";
    when 16#1496# => romdata <= X"88092003";
    when 16#1497# => romdata <= X"8736A012";
    when 16#1498# => romdata <= X"88113FF8";
    when 16#1499# => romdata <= X"8608E03F";
    when 16#149A# => romdata <= X"8536A00C";
    when 16#149B# => romdata <= X"8610FF80";
    when 16#149C# => romdata <= X"8408A03F";
    when 16#149D# => romdata <= X"820EAFC0";
    when 16#149E# => romdata <= X"8410BF80";
    when 16#149F# => romdata <= X"83386006";
    when 16#14A0# => romdata <= X"82107F80";
    when 16#14A1# => romdata <= X"DA2E6004";
    when 16#14A2# => romdata <= X"C82E4000";
    when 16#14A3# => romdata <= X"C62E6001";
    when 16#14A4# => romdata <= X"C42E6002";
    when 16#14A5# => romdata <= X"C22E6003";
    when 16#14A6# => romdata <= X"81C7E008";
    when 16#14A7# => romdata <= X"91E82005";
    when 16#14A8# => romdata <= X"8608E0FF";
    when 16#14A9# => romdata <= X"80A0E00F";
    when 16#14AA# => romdata <= X"38800050";
    when 16#14AB# => romdata <= X"8200607F";
    when 16#14AC# => romdata <= X"8206BF80";
    when 16#14AD# => romdata <= X"820860FF";
    when 16#14AE# => romdata <= X"80A0607C";
    when 16#14AF# => romdata <= X"08800007";
    when 16#14B0# => romdata <= X"8210001A";
    when 16#14B1# => romdata <= X"8606BFC0";
    when 16#14B2# => romdata <= X"8608E0FF";
    when 16#14B3# => romdata <= X"80A0E03E";
    when 16#14B4# => romdata <= X"38800033";
    when 16#14B5# => romdata <= X"B0103FFF";
    when 16#14B6# => romdata <= X"C22E6001";
    when 16#14B7# => romdata <= X"C42E4000";
    when 16#14B8# => romdata <= X"81C7E008";
    when 16#14B9# => romdata <= X"91E82002";
    when 16#14BA# => romdata <= X"90142120";
    when 16#14BB# => romdata <= X"13100032";
    when 16#14BC# => romdata <= X"7FFFF4B1";
    when 16#14BD# => romdata <= X"92126098";
    when 16#14BE# => romdata <= X"80A22000";
    when 16#14BF# => romdata <= X"1280000E";
    when 16#14C0# => romdata <= X"80A66000";
    when 16#14C1# => romdata <= X"02BFFFAE";
    when 16#14C2# => romdata <= X"833EA008";
    when 16#14C3# => romdata <= X"808860FF";
    when 16#14C4# => romdata <= X"22BFFFA6";
    when 16#14C5# => romdata <= X"F42E4000";
    when 16#14C6# => romdata <= X"8400605F";
    when 16#14C7# => romdata <= X"8408A0FF";
    when 16#14C8# => romdata <= X"80A0A05D";
    when 16#14C9# => romdata <= X"0880006C";
    when 16#14CA# => romdata <= X"8406A05F";
    when 16#14CB# => romdata <= X"81C7E008";
    when 16#14CC# => romdata <= X"91E83FFF";
    when 16#14CD# => romdata <= X"90142120";
    when 16#14CE# => romdata <= X"13100032";
    when 16#14CF# => romdata <= X"7FFFF49E";
    when 16#14D0# => romdata <= X"921260A0";
    when 16#14D1# => romdata <= X"80A22000";
    when 16#14D2# => romdata <= X"12BFFF9B";
    when 16#14D3# => romdata <= X"80A66000";
    when 16#14D4# => romdata <= X"02800013";
    when 16#14D5# => romdata <= X"B0102001";
    when 16#14D6# => romdata <= X"833EA008";
    when 16#14D7# => romdata <= X"868860FF";
    when 16#14D8# => romdata <= X"12800041";
    when 16#14D9# => romdata <= X"8410001A";
    when 16#14DA# => romdata <= X"C206C000";
    when 16#14DB# => romdata <= X"80A06000";
    when 16#14DC# => romdata <= X"0280000A";
    when 16#14DD# => romdata <= X"8210201B";
    when 16#14DE# => romdata <= X"C026C000";
    when 16#14DF# => romdata <= X"C22E4000";
    when 16#14E0# => romdata <= X"82102028";
    when 16#14E1# => romdata <= X"B0102004";
    when 16#14E2# => romdata <= X"C22E6001";
    when 16#14E3# => romdata <= X"82102042";
    when 16#14E4# => romdata <= X"C22E6002";
    when 16#14E5# => romdata <= X"B2066003";
    when 16#14E6# => romdata <= X"C42E4000";
    when 16#14E7# => romdata <= X"81C7E008";
    when 16#14E8# => romdata <= X"81E80000";
    when 16#14E9# => romdata <= X"033FFFCA";
    when 16#14EA# => romdata <= X"82068001";
    when 16#14EB# => romdata <= X"80A067FF";
    when 16#14EC# => romdata <= X"08BFFFDF";
    when 16#14ED# => romdata <= X"860EA03F";
    when 16#14EE# => romdata <= X"8536A00C";
    when 16#14EF# => romdata <= X"8610FF80";
    when 16#14F0# => romdata <= X"8408A00F";
    when 16#14F1# => romdata <= X"820EAFC0";
    when 16#14F2# => romdata <= X"8410BFE0";
    when 16#14F3# => romdata <= X"83386006";
    when 16#14F4# => romdata <= X"82107F80";
    when 16#14F5# => romdata <= X"C62E6002";
    when 16#14F6# => romdata <= X"C42E4000";
    when 16#14F7# => romdata <= X"C22E6001";
    when 16#14F8# => romdata <= X"81C7E008";
    when 16#14F9# => romdata <= X"91E82003";
    when 16#14FA# => romdata <= X"820860FF";
    when 16#14FB# => romdata <= X"80A0601E";
    when 16#14FC# => romdata <= X"08BFFFB1";
    when 16#14FD# => romdata <= X"8206BF80";
    when 16#14FE# => romdata <= X"81C7E008";
    when 16#14FF# => romdata <= X"91E83FFF";
    when 16#1500# => romdata <= X"980EA03F";
    when 16#1501# => romdata <= X"9B36A01E";
    when 16#1502# => romdata <= X"98133F80";
    when 16#1503# => romdata <= X"9A0B6001";
    when 16#1504# => romdata <= X"8936A018";
    when 16#1505# => romdata <= X"9A137FFC";
    when 16#1506# => romdata <= X"8809203F";
    when 16#1507# => romdata <= X"8736A012";
    when 16#1508# => romdata <= X"88113F80";
    when 16#1509# => romdata <= X"8608E03F";
    when 16#150A# => romdata <= X"8536A00C";
    when 16#150B# => romdata <= X"8610FF80";
    when 16#150C# => romdata <= X"8408A03F";
    when 16#150D# => romdata <= X"820EAFC0";
    when 16#150E# => romdata <= X"8410BF80";
    when 16#150F# => romdata <= X"83386006";
    when 16#1510# => romdata <= X"82107F80";
    when 16#1511# => romdata <= X"D82E6005";
    when 16#1512# => romdata <= X"DA2E4000";
    when 16#1513# => romdata <= X"C82E6001";
    when 16#1514# => romdata <= X"C62E6002";
    when 16#1515# => romdata <= X"C42E6003";
    when 16#1516# => romdata <= X"C22E6004";
    when 16#1517# => romdata <= X"81C7E008";
    when 16#1518# => romdata <= X"91E82006";
    when 16#1519# => romdata <= X"82007FDF";
    when 16#151A# => romdata <= X"820860FF";
    when 16#151B# => romdata <= X"80A0605D";
    when 16#151C# => romdata <= X"18BFFFCB";
    when 16#151D# => romdata <= X"B0103FFF";
    when 16#151E# => romdata <= X"8206BFDF";
    when 16#151F# => romdata <= X"820860FF";
    when 16#1520# => romdata <= X"80A0605D";
    when 16#1521# => romdata <= X"18800012";
    when 16#1522# => romdata <= X"01000000";
    when 16#1523# => romdata <= X"C206C000";
    when 16#1524# => romdata <= X"80A06000";
    when 16#1525# => romdata <= X"1280000C";
    when 16#1526# => romdata <= X"B0102002";
    when 16#1527# => romdata <= X"82102001";
    when 16#1528# => romdata <= X"C226C000";
    when 16#1529# => romdata <= X"8210201B";
    when 16#152A# => romdata <= X"C22E4000";
    when 16#152B# => romdata <= X"82102024";
    when 16#152C# => romdata <= X"B0102005";
    when 16#152D# => romdata <= X"C22E6001";
    when 16#152E# => romdata <= X"82102042";
    when 16#152F# => romdata <= X"C22E6002";
    when 16#1530# => romdata <= X"B2066003";
    when 16#1531# => romdata <= X"C42E6001";
    when 16#1532# => romdata <= X"C62E4000";
    when 16#1533# => romdata <= X"81C7E008";
    when 16#1534# => romdata <= X"81E80000";
    when 16#1535# => romdata <= X"8408A0FF";
    when 16#1536# => romdata <= X"80A0A05D";
    when 16#1537# => romdata <= X"38BFFFB0";
    when 16#1538# => romdata <= X"B0103FFF";
    when 16#1539# => romdata <= X"F42E6001";
    when 16#153A# => romdata <= X"C22E4000";
    when 16#153B# => romdata <= X"81C7E008";
    when 16#153C# => romdata <= X"91E82002";
    when 16#153D# => romdata <= X"9DE3BFA0";
    when 16#153E# => romdata <= X"23100032";
    when 16#153F# => romdata <= X"D00462C8";
    when 16#1540# => romdata <= X"80A22000";
    when 16#1541# => romdata <= X"02800006";
    when 16#1542# => romdata <= X"A0100018";
    when 16#1543# => romdata <= X"C2022038";
    when 16#1544# => romdata <= X"80A06000";
    when 16#1545# => romdata <= X"02800020";
    when 16#1546# => romdata <= X"01000000";
    when 16#1547# => romdata <= X"C214200C";
    when 16#1548# => romdata <= X"85286010";
    when 16#1549# => romdata <= X"8530A010";
    when 16#154A# => romdata <= X"8088A008";
    when 16#154B# => romdata <= X"02800022";
    when 16#154C# => romdata <= X"86100001";
    when 16#154D# => romdata <= X"C4042010";
    when 16#154E# => romdata <= X"80A0A000";
    when 16#154F# => romdata <= X"0280001A";
    when 16#1550# => romdata <= X"01000000";
    when 16#1551# => romdata <= X"C214200C";
    when 16#1552# => romdata <= X"80886001";
    when 16#1553# => romdata <= X"1280000C";
    when 16#1554# => romdata <= X"80886002";
    when 16#1555# => romdata <= X"02800006";
    when 16#1556# => romdata <= X"82102000";
    when 16#1557# => romdata <= X"C2242008";
    when 16#1558# => romdata <= X"B0102000";
    when 16#1559# => romdata <= X"81C7E008";
    when 16#155A# => romdata <= X"81E80000";
    when 16#155B# => romdata <= X"C2042014";
    when 16#155C# => romdata <= X"C2242008";
    when 16#155D# => romdata <= X"81C7E008";
    when 16#155E# => romdata <= X"91E82000";
    when 16#155F# => romdata <= X"C2042014";
    when 16#1560# => romdata <= X"82200001";
    when 16#1561# => romdata <= X"C0242008";
    when 16#1562# => romdata <= X"C2242018";
    when 16#1563# => romdata <= X"81C7E008";
    when 16#1564# => romdata <= X"91E82000";
    when 16#1565# => romdata <= X"40000621";
    when 16#1566# => romdata <= X"01000000";
    when 16#1567# => romdata <= X"10BFFFE1";
    when 16#1568# => romdata <= X"C214200C";
    when 16#1569# => romdata <= X"4000091A";
    when 16#156A# => romdata <= X"90100010";
    when 16#156B# => romdata <= X"10BFFFE7";
    when 16#156C# => romdata <= X"C214200C";
    when 16#156D# => romdata <= X"8088A010";
    when 16#156E# => romdata <= X"02BFFFEB";
    when 16#156F# => romdata <= X"B0103FFF";
    when 16#1570# => romdata <= X"8088A004";
    when 16#1571# => romdata <= X"32800006";
    when 16#1572# => romdata <= X"D2042030";
    when 16#1573# => romdata <= X"8610E008";
    when 16#1574# => romdata <= X"C4042010";
    when 16#1575# => romdata <= X"10BFFFD9";
    when 16#1576# => romdata <= X"C634200C";
    when 16#1577# => romdata <= X"80A26000";
    when 16#1578# => romdata <= X"0280000B";
    when 16#1579# => romdata <= X"86087FDB";
    when 16#157A# => romdata <= X"84042040";
    when 16#157B# => romdata <= X"80A24002";
    when 16#157C# => romdata <= X"22800007";
    when 16#157D# => romdata <= X"C0242030";
    when 16#157E# => romdata <= X"400006B9";
    when 16#157F# => romdata <= X"D00462C8";
    when 16#1580# => romdata <= X"C214200C";
    when 16#1581# => romdata <= X"C0242030";
    when 16#1582# => romdata <= X"86087FDB";
    when 16#1583# => romdata <= X"C4042010";
    when 16#1584# => romdata <= X"C0242004";
    when 16#1585# => romdata <= X"C634200C";
    when 16#1586# => romdata <= X"8610E008";
    when 16#1587# => romdata <= X"C4240000";
    when 16#1588# => romdata <= X"10BFFFC6";
    when 16#1589# => romdata <= X"C634200C";
    when 16#158A# => romdata <= X"9DE3BFA0";
    when 16#158B# => romdata <= X"C2062010";
    when 16#158C# => romdata <= X"E6066010";
    when 16#158D# => romdata <= X"A0100018";
    when 16#158E# => romdata <= X"80A4C001";
    when 16#158F# => romdata <= X"1480007F";
    when 16#1590# => romdata <= X"B0102000";
    when 16#1591# => romdata <= X"BA04E003";
    when 16#1592# => romdata <= X"BB2F6002";
    when 16#1593# => romdata <= X"8204001D";
    when 16#1594# => romdata <= X"BA06401D";
    when 16#1595# => romdata <= X"F4006004";
    when 16#1596# => romdata <= X"D2076004";
    when 16#1597# => romdata <= X"92026001";
    when 16#1598# => romdata <= X"9010001A";
    when 16#1599# => romdata <= X"4000112F";
    when 16#159A# => romdata <= X"A604FFFF";
    when 16#159B# => romdata <= X"BA076004";
    when 16#159C# => romdata <= X"B0922000";
    when 16#159D# => romdata <= X"A2066014";
    when 16#159E# => romdata <= X"0280003B";
    when 16#159F# => romdata <= X"B8042014";
    when 16#15A0# => romdata <= X"2B00003F";
    when 16#15A1# => romdata <= X"A8100011";
    when 16#15A2# => romdata <= X"AA1563FF";
    when 16#15A3# => romdata <= X"A410001C";
    when 16#15A4# => romdata <= X"AC102000";
    when 16#15A5# => romdata <= X"B6102000";
    when 16#15A6# => romdata <= X"EE050000";
    when 16#15A7# => romdata <= X"920DC015";
    when 16#15A8# => romdata <= X"400010E6";
    when 16#15A9# => romdata <= X"90100018";
    when 16#15AA# => romdata <= X"9335E010";
    when 16#15AB# => romdata <= X"AC058008";
    when 16#15AC# => romdata <= X"400010E2";
    when 16#15AD# => romdata <= X"90100018";
    when 16#15AE# => romdata <= X"C2048000";
    when 16#15AF# => romdata <= X"87306010";
    when 16#15B0# => romdata <= X"82084015";
    when 16#15B1# => romdata <= X"B606C001";
    when 16#15B2# => romdata <= X"840D8015";
    when 16#15B3# => romdata <= X"AD35A010";
    when 16#15B4# => romdata <= X"8426C002";
    when 16#15B5# => romdata <= X"AC058008";
    when 16#15B6# => romdata <= X"8338A010";
    when 16#15B7# => romdata <= X"880D8015";
    when 16#15B8# => romdata <= X"8620C004";
    when 16#15B9# => romdata <= X"B600C001";
    when 16#15BA# => romdata <= X"C434A002";
    when 16#15BB# => romdata <= X"A8052004";
    when 16#15BC# => romdata <= X"F6348000";
    when 16#15BD# => romdata <= X"80A74014";
    when 16#15BE# => romdata <= X"A404A004";
    when 16#15BF# => romdata <= X"AD35A010";
    when 16#15C0# => romdata <= X"1ABFFFE6";
    when 16#15C1# => romdata <= X"B73EE010";
    when 16#15C2# => romdata <= X"80A6A000";
    when 16#15C3# => romdata <= X"12800017";
    when 16#15C4# => romdata <= X"92100019";
    when 16#15C5# => romdata <= X"8404E004";
    when 16#15C6# => romdata <= X"8528A002";
    when 16#15C7# => romdata <= X"82040002";
    when 16#15C8# => romdata <= X"80A70001";
    when 16#15C9# => romdata <= X"3A800011";
    when 16#15CA# => romdata <= X"E6242010";
    when 16#15CB# => romdata <= X"C4040002";
    when 16#15CC# => romdata <= X"80A0A000";
    when 16#15CD# => romdata <= X"02800008";
    when 16#15CE# => romdata <= X"82007FFC";
    when 16#15CF# => romdata <= X"1080000B";
    when 16#15D0# => romdata <= X"E6242010";
    when 16#15D1# => romdata <= X"C4004000";
    when 16#15D2# => romdata <= X"80A0A000";
    when 16#15D3# => romdata <= X"12800005";
    when 16#15D4# => romdata <= X"82007FFC";
    when 16#15D5# => romdata <= X"80A70001";
    when 16#15D6# => romdata <= X"0ABFFFFB";
    when 16#15D7# => romdata <= X"A604FFFF";
    when 16#15D8# => romdata <= X"E6242010";
    when 16#15D9# => romdata <= X"92100019";
    when 16#15DA# => romdata <= X"40000A6C";
    when 16#15DB# => romdata <= X"90100010";
    when 16#15DC# => romdata <= X"80A22000";
    when 16#15DD# => romdata <= X"06800031";
    when 16#15DE# => romdata <= X"1700003F";
    when 16#15DF# => romdata <= X"B0062001";
    when 16#15E0# => romdata <= X"9612E3FF";
    when 16#15E1# => romdata <= X"8210001C";
    when 16#15E2# => romdata <= X"98102000";
    when 16#15E3# => romdata <= X"C8044000";
    when 16#15E4# => romdata <= X"DA004000";
    when 16#15E5# => romdata <= X"87336010";
    when 16#15E6# => romdata <= X"85312010";
    when 16#15E7# => romdata <= X"8809000B";
    when 16#15E8# => romdata <= X"8420C002";
    when 16#15E9# => romdata <= X"860B400B";
    when 16#15EA# => romdata <= X"8620C004";
    when 16#15EB# => romdata <= X"8600C00C";
    when 16#15EC# => romdata <= X"8938E010";
    when 16#15ED# => romdata <= X"84008004";
    when 16#15EE# => romdata <= X"C6306002";
    when 16#15EF# => romdata <= X"A2046004";
    when 16#15F0# => romdata <= X"C4304000";
    when 16#15F1# => romdata <= X"80A74011";
    when 16#15F2# => romdata <= X"82006004";
    when 16#15F3# => romdata <= X"1ABFFFF0";
    when 16#15F4# => romdata <= X"9938A010";
    when 16#15F5# => romdata <= X"8404E004";
    when 16#15F6# => romdata <= X"8528A002";
    when 16#15F7# => romdata <= X"82040002";
    when 16#15F8# => romdata <= X"C6006004";
    when 16#15F9# => romdata <= X"80A0E000";
    when 16#15FA# => romdata <= X"12800014";
    when 16#15FB# => romdata <= X"80A70001";
    when 16#15FC# => romdata <= X"3A800012";
    when 16#15FD# => romdata <= X"E6242010";
    when 16#15FE# => romdata <= X"C4040002";
    when 16#15FF# => romdata <= X"80A0A000";
    when 16#1600# => romdata <= X"2280000A";
    when 16#1601# => romdata <= X"82007FFC";
    when 16#1602# => romdata <= X"E6242010";
    when 16#1603# => romdata <= X"81C7E008";
    when 16#1604# => romdata <= X"81E80000";
    when 16#1605# => romdata <= X"C4004000";
    when 16#1606# => romdata <= X"80A0A000";
    when 16#1607# => romdata <= X"32800007";
    when 16#1608# => romdata <= X"E6242010";
    when 16#1609# => romdata <= X"82007FFC";
    when 16#160A# => romdata <= X"80A70001";
    when 16#160B# => romdata <= X"0ABFFFFA";
    when 16#160C# => romdata <= X"A604FFFF";
    when 16#160D# => romdata <= X"E6242010";
    when 16#160E# => romdata <= X"81C7E008";
    when 16#160F# => romdata <= X"81E80000";
    when 16#1610# => romdata <= X"9DE3BF60";
    when 16#1611# => romdata <= X"C2062040";
    when 16#1612# => romdata <= X"F227BFC8";
    when 16#1613# => romdata <= X"F427BFCC";
    when 16#1614# => romdata <= X"80A06000";
    when 16#1615# => romdata <= X"E207A05C";
    when 16#1616# => romdata <= X"E007A060";
    when 16#1617# => romdata <= X"02800010";
    when 16#1618# => romdata <= X"D11FBFC8";
    when 16#1619# => romdata <= X"C4062044";
    when 16#161A# => romdata <= X"C4206004";
    when 16#161B# => romdata <= X"86102001";
    when 16#161C# => romdata <= X"D127BFD4";
    when 16#161D# => romdata <= X"C4062044";
    when 16#161E# => romdata <= X"8528C002";
    when 16#161F# => romdata <= X"C4206008";
    when 16#1620# => romdata <= X"D327BFD0";
    when 16#1621# => romdata <= X"92100001";
    when 16#1622# => romdata <= X"400009BF";
    when 16#1623# => romdata <= X"90100018";
    when 16#1624# => romdata <= X"D307BFD0";
    when 16#1625# => romdata <= X"C0262040";
    when 16#1626# => romdata <= X"D107BFD4";
    when 16#1627# => romdata <= X"D127BFC4";
    when 16#1628# => romdata <= X"E407BFC4";
    when 16#1629# => romdata <= X"80A4A000";
    when 16#162A# => romdata <= X"0680003E";
    when 16#162B# => romdata <= X"82102001";
    when 16#162C# => romdata <= X"C0244000";
    when 16#162D# => romdata <= X"031FFC00";
    when 16#162E# => romdata <= X"840C8001";
    when 16#162F# => romdata <= X"80A08001";
    when 16#1630# => romdata <= X"02800023";
    when 16#1631# => romdata <= X"23100032";
    when 16#1632# => romdata <= X"95A00028";
    when 16#1633# => romdata <= X"D91C6060";
    when 16#1634# => romdata <= X"97A00029";
    when 16#1635# => romdata <= X"81AA8A4C";
    when 16#1636# => romdata <= X"01000000";
    when 16#1637# => romdata <= X"03800037";
    when 16#1638# => romdata <= X"82102001";
    when 16#1639# => romdata <= X"C2274000";
    when 16#163A# => romdata <= X"31100032";
    when 16#163B# => romdata <= X"80A42000";
    when 16#163C# => romdata <= X"02800015";
    when 16#163D# => romdata <= X"B0162048";
    when 16#163E# => romdata <= X"31100032";
    when 16#163F# => romdata <= X"B0162049";
    when 16#1640# => romdata <= X"F0240000";
    when 16#1641# => romdata <= X"81C7E008";
    when 16#1642# => romdata <= X"91EE3FFF";
    when 16#1643# => romdata <= X"8400A001";
    when 16#1644# => romdata <= X"C4284000";
    when 16#1645# => romdata <= X"E627BFEC";
    when 16#1646# => romdata <= X"90100018";
    when 16#1647# => romdata <= X"4000099A";
    when 16#1648# => romdata <= X"92100014";
    when 16#1649# => romdata <= X"C02C8000";
    when 16#164A# => romdata <= X"80A42000";
    when 16#164B# => romdata <= X"B0100015";
    when 16#164C# => romdata <= X"C407BFEC";
    when 16#164D# => romdata <= X"8200A001";
    when 16#164E# => romdata <= X"02800003";
    when 16#164F# => romdata <= X"C2274000";
    when 16#1650# => romdata <= X"E4240000";
    when 16#1651# => romdata <= X"81C7E008";
    when 16#1652# => romdata <= X"81E80000";
    when 16#1653# => romdata <= X"D327BFC4";
    when 16#1654# => romdata <= X"03000009";
    when 16#1655# => romdata <= X"8210630F";
    when 16#1656# => romdata <= X"C2274000";
    when 16#1657# => romdata <= X"C407BFC4";
    when 16#1658# => romdata <= X"80A0A000";
    when 16#1659# => romdata <= X"028000FA";
    when 16#165A# => romdata <= X"033FFC00";
    when 16#165B# => romdata <= X"31100032";
    when 16#165C# => romdata <= X"B0162040";
    when 16#165D# => romdata <= X"80A42000";
    when 16#165E# => romdata <= X"02800008";
    when 16#165F# => romdata <= X"01000000";
    when 16#1660# => romdata <= X"C24E2003";
    when 16#1661# => romdata <= X"80A06000";
    when 16#1662# => romdata <= X"02800003";
    when 16#1663# => romdata <= X"82062003";
    when 16#1664# => romdata <= X"82062008";
    when 16#1665# => romdata <= X"C2240000";
    when 16#1666# => romdata <= X"81C7E008";
    when 16#1667# => romdata <= X"81E80000";
    when 16#1668# => romdata <= X"C2244000";
    when 16#1669# => romdata <= X"03200000";
    when 16#166A# => romdata <= X"A42C8001";
    when 16#166B# => romdata <= X"E427BFC4";
    when 16#166C# => romdata <= X"10BFFFC1";
    when 16#166D# => romdata <= X"D107BFC4";
    when 16#166E# => romdata <= X"D53FBFC8";
    when 16#166F# => romdata <= X"D127BFD4";
    when 16#1670# => romdata <= X"D327BFD0";
    when 16#1671# => romdata <= X"D127BFDC";
    when 16#1672# => romdata <= X"D327BFD8";
    when 16#1673# => romdata <= X"90100018";
    when 16#1674# => romdata <= X"9607BFF8";
    when 16#1675# => romdata <= X"D81FBFC8";
    when 16#1676# => romdata <= X"9210000C";
    when 16#1677# => romdata <= X"9410000D";
    when 16#1678# => romdata <= X"40000ABB";
    when 16#1679# => romdata <= X"9807BFFC";
    when 16#167A# => romdata <= X"8934A014";
    when 16#167B# => romdata <= X"A8100008";
    when 16#167C# => romdata <= X"888927FF";
    when 16#167D# => romdata <= X"D107BFD4";
    when 16#167E# => romdata <= X"D307BFD0";
    when 16#167F# => romdata <= X"D507BFDC";
    when 16#1680# => romdata <= X"128000D9";
    when 16#1681# => romdata <= X"D707BFD8";
    when 16#1682# => romdata <= X"D327BFC4";
    when 16#1683# => romdata <= X"C207BFFC";
    when 16#1684# => romdata <= X"C607BFF8";
    when 16#1685# => romdata <= X"86004003";
    when 16#1686# => romdata <= X"8800E432";
    when 16#1687# => romdata <= X"84200004";
    when 16#1688# => romdata <= X"80A12020";
    when 16#1689# => romdata <= X"DA07BFC4";
    when 16#168A# => romdata <= X"04800007";
    when 16#168B# => romdata <= X"852B4002";
    when 16#168C# => romdata <= X"8600E412";
    when 16#168D# => romdata <= X"84200004";
    when 16#168E# => romdata <= X"87334003";
    when 16#168F# => romdata <= X"852C8002";
    when 16#1690# => romdata <= X"84108003";
    when 16#1691# => romdata <= X"C427BFC4";
    when 16#1692# => romdata <= X"80A0A000";
    when 16#1693# => romdata <= X"DD07BFC4";
    when 16#1694# => romdata <= X"06800369";
    when 16#1695# => romdata <= X"99A0190E";
    when 16#1696# => romdata <= X"D93FBFC8";
    when 16#1697# => romdata <= X"88013BCD";
    when 16#1698# => romdata <= X"D81FBFC8";
    when 16#1699# => romdata <= X"8610000D";
    when 16#169A# => romdata <= X"1B3F8400";
    when 16#169B# => romdata <= X"8410000C";
    when 16#169C# => romdata <= X"84034002";
    when 16#169D# => romdata <= X"9A102001";
    when 16#169E# => romdata <= X"DA27BFE8";
    when 16#169F# => romdata <= X"C43FBFC8";
    when 16#16A0# => romdata <= X"C827BFC4";
    when 16#16A1# => romdata <= X"1B100032";
    when 16#16A2# => romdata <= X"DD1B60C0";
    when 16#16A3# => romdata <= X"05100032";
    when 16#16A4# => romdata <= X"D91FBFC8";
    when 16#16A5# => romdata <= X"9DA308CE";
    when 16#16A6# => romdata <= X"D918A0C8";
    when 16#16A7# => romdata <= X"9DA3894C";
    when 16#16A8# => romdata <= X"DB07BFC4";
    when 16#16A9# => romdata <= X"A1A0190D";
    when 16#16AA# => romdata <= X"05100032";
    when 16#16AB# => romdata <= X"D918A0D0";
    when 16#16AC# => romdata <= X"9DA3884C";
    when 16#16AD# => romdata <= X"05100032";
    when 16#16AE# => romdata <= X"D918A0D8";
    when 16#16AF# => romdata <= X"99A4094C";
    when 16#16B0# => romdata <= X"99A3884C";
    when 16#16B1# => romdata <= X"DD1C6060";
    when 16#16B2# => romdata <= X"81AB0ACE";
    when 16#16B3# => romdata <= X"9DA01A4C";
    when 16#16B4# => romdata <= X"DD27BFC4";
    when 16#16B5# => romdata <= X"01000000";
    when 16#16B6# => romdata <= X"19800007";
    when 16#16B7# => romdata <= X"E607BFC4";
    when 16#16B8# => romdata <= X"9DA0190E";
    when 16#16B9# => romdata <= X"81AB8A4C";
    when 16#16BA# => romdata <= X"01000000";
    when 16#16BB# => romdata <= X"23800002";
    when 16#16BC# => romdata <= X"A604FFFF";
    when 16#16BD# => romdata <= X"84102001";
    when 16#16BE# => romdata <= X"80A4E016";
    when 16#16BF# => romdata <= X"1880000B";
    when 16#16C0# => romdata <= X"C427BFF4";
    when 16#16C1# => romdata <= X"852CE003";
    when 16#16C2# => romdata <= X"07100032";
    when 16#16C3# => romdata <= X"8610E150";
    when 16#16C4# => romdata <= X"D918C002";
    when 16#16C5# => romdata <= X"81AA8ACC";
    when 16#16C6# => romdata <= X"01000000";
    when 16#16C7# => romdata <= X"19800003";
    when 16#16C8# => romdata <= X"C027BFF4";
    when 16#16C9# => romdata <= X"A604FFFF";
    when 16#16CA# => romdata <= X"82007FFF";
    when 16#16CB# => romdata <= X"B4102000";
    when 16#16CC# => romdata <= X"82204004";
    when 16#16CD# => romdata <= X"80A06000";
    when 16#16CE# => romdata <= X"06800004";
    when 16#16CF# => romdata <= X"B2200001";
    when 16#16D0# => romdata <= X"B4100001";
    when 16#16D1# => romdata <= X"B2102000";
    when 16#16D2# => romdata <= X"80A4E000";
    when 16#16D3# => romdata <= X"068001D9";
    when 16#16D4# => romdata <= X"86200013";
    when 16#16D5# => romdata <= X"E627BFE4";
    when 16#16D6# => romdata <= X"C027BFF0";
    when 16#16D7# => romdata <= X"B4068013";
    when 16#16D8# => romdata <= X"80A6E009";
    when 16#16D9# => romdata <= X"1880008C";
    when 16#16DA# => romdata <= X"86103FFF";
    when 16#16DB# => romdata <= X"80A6E005";
    when 16#16DC# => romdata <= X"04800004";
    when 16#16DD# => romdata <= X"A4102001";
    when 16#16DE# => romdata <= X"B606FFFC";
    when 16#16DF# => romdata <= X"A4102000";
    when 16#16E0# => romdata <= X"80A6E003";
    when 16#16E1# => romdata <= X"0280000A";
    when 16#16E2# => romdata <= X"AE102000";
    when 16#16E3# => romdata <= X"048001D3";
    when 16#16E4# => romdata <= X"80A6E002";
    when 16#16E5# => romdata <= X"80A6E004";
    when 16#16E6# => romdata <= X"0280031B";
    when 16#16E7# => romdata <= X"80A6E005";
    when 16#16E8# => romdata <= X"128001D0";
    when 16#16E9# => romdata <= X"88103FFF";
    when 16#16EA# => romdata <= X"AE102001";
    when 16#16EB# => romdata <= X"9A04C01C";
    when 16#16EC# => romdata <= X"88036001";
    when 16#16ED# => romdata <= X"AC912000";
    when 16#16EE# => romdata <= X"04800348";
    when 16#16EF# => romdata <= X"DA27BFE0";
    when 16#16F0# => romdata <= X"C0262044";
    when 16#16F1# => romdata <= X"80A12017";
    when 16#16F2# => romdata <= X"84102001";
    when 16#16F3# => romdata <= X"088003D5";
    when 16#16F4# => romdata <= X"82102004";
    when 16#16F5# => romdata <= X"92100002";
    when 16#16F6# => romdata <= X"83286001";
    when 16#16F7# => romdata <= X"86006014";
    when 16#16F8# => romdata <= X"80A0C004";
    when 16#16F9# => romdata <= X"08BFFFFC";
    when 16#16FA# => romdata <= X"8400A001";
    when 16#16FB# => romdata <= X"80A5A00F";
    when 16#16FC# => romdata <= X"D2262044";
    when 16#16FD# => romdata <= X"82402000";
    when 16#16FE# => romdata <= X"D127BFD4";
    when 16#16FF# => romdata <= X"A4084012";
    when 16#1700# => romdata <= X"D327BFD0";
    when 16#1701# => romdata <= X"D527BFDC";
    when 16#1702# => romdata <= X"D727BFD8";
    when 16#1703# => romdata <= X"40000A06";
    when 16#1704# => romdata <= X"90100018";
    when 16#1705# => romdata <= X"D0262040";
    when 16#1706# => romdata <= X"AA100008";
    when 16#1707# => romdata <= X"808CA0FF";
    when 16#1708# => romdata <= X"D107BFD4";
    when 16#1709# => romdata <= X"D307BFD0";
    when 16#170A# => romdata <= X"D507BFDC";
    when 16#170B# => romdata <= X"12800070";
    when 16#170C# => romdata <= X"D707BFD8";
    when 16#170D# => romdata <= X"80A4E00E";
    when 16#170E# => romdata <= X"148000CC";
    when 16#170F# => romdata <= X"C207BFF8";
    when 16#1710# => romdata <= X"80A06000";
    when 16#1711# => romdata <= X"068000C9";
    when 16#1712# => romdata <= X"05100032";
    when 16#1713# => romdata <= X"832CE003";
    when 16#1714# => romdata <= X"80A5A000";
    when 16#1715# => romdata <= X"8410A150";
    when 16#1716# => romdata <= X"0480026D";
    when 16#1717# => romdata <= X"D9188001";
    when 16#1718# => romdata <= X"95A209CC";
    when 16#1719# => romdata <= X"80A5A001";
    when 16#171A# => romdata <= X"A4056001";
    when 16#171B# => romdata <= X"95A01A4A";
    when 16#171C# => romdata <= X"D527BFC4";
    when 16#171D# => romdata <= X"9DA0190A";
    when 16#171E# => romdata <= X"9DA3894C";
    when 16#171F# => romdata <= X"91A208CE";
    when 16#1720# => romdata <= X"D807BFC4";
    when 16#1721# => romdata <= X"82032030";
    when 16#1722# => romdata <= X"02800021";
    when 16#1723# => romdata <= X"C22D4000";
    when 16#1724# => romdata <= X"1B100032";
    when 16#1725# => romdata <= X"D51B60E8";
    when 16#1726# => romdata <= X"91A2094A";
    when 16#1727# => romdata <= X"D51C6060";
    when 16#1728# => romdata <= X"81AA0A4A";
    when 16#1729# => romdata <= X"01000000";
    when 16#172A# => romdata <= X"13800027";
    when 16#172B# => romdata <= X"82102001";
    when 16#172C# => romdata <= X"861360E8";
    when 16#172D# => romdata <= X"10800009";
    when 16#172E# => romdata <= X"A2146060";
    when 16#172F# => romdata <= X"D518C000";
    when 16#1730# => romdata <= X"91A2094A";
    when 16#1731# => romdata <= X"D51C4000";
    when 16#1732# => romdata <= X"81AA0A4A";
    when 16#1733# => romdata <= X"01000000";
    when 16#1734# => romdata <= X"33BFFF12";
    when 16#1735# => romdata <= X"E627BFEC";
    when 16#1736# => romdata <= X"95A209CC";
    when 16#1737# => romdata <= X"82006001";
    when 16#1738# => romdata <= X"80A58001";
    when 16#1739# => romdata <= X"95A01A4A";
    when 16#173A# => romdata <= X"D527BFC4";
    when 16#173B# => romdata <= X"9DA0190A";
    when 16#173C# => romdata <= X"9DA3894C";
    when 16#173D# => romdata <= X"91A208CE";
    when 16#173E# => romdata <= X"C807BFC4";
    when 16#173F# => romdata <= X"84012030";
    when 16#1740# => romdata <= X"C42C8000";
    when 16#1741# => romdata <= X"12BFFFEE";
    when 16#1742# => romdata <= X"A404A001";
    when 16#1743# => romdata <= X"91A20848";
    when 16#1744# => romdata <= X"81AB0AC8";
    when 16#1745# => romdata <= X"01000000";
    when 16#1746# => romdata <= X"29800226";
    when 16#1747# => romdata <= X"C24CBFFF";
    when 16#1748# => romdata <= X"81AB0A48";
    when 16#1749# => romdata <= X"01000000";
    when 16#174A# => romdata <= X"23BFFEFC";
    when 16#174B# => romdata <= X"E627BFEC";
    when 16#174C# => romdata <= X"D527BFC4";
    when 16#174D# => romdata <= X"DA07BFC4";
    when 16#174E# => romdata <= X"808B6001";
    when 16#174F# => romdata <= X"3280021D";
    when 16#1750# => romdata <= X"C24CBFFF";
    when 16#1751# => romdata <= X"10BFFEF5";
    when 16#1752# => romdata <= X"E627BFEC";
    when 16#1753# => romdata <= X"31100032";
    when 16#1754# => romdata <= X"80AC8001";
    when 16#1755# => romdata <= X"02BFFF08";
    when 16#1756# => romdata <= X"B01620A8";
    when 16#1757# => romdata <= X"10BFFF05";
    when 16#1758# => romdata <= X"31100032";
    when 16#1759# => romdata <= X"D53FBFC8";
    when 16#175A# => romdata <= X"030FFC00";
    when 16#175B# => romdata <= X"88013C01";
    when 16#175C# => romdata <= X"C027BFE8";
    when 16#175D# => romdata <= X"D81FBFC8";
    when 16#175E# => romdata <= X"8410000C";
    when 16#175F# => romdata <= X"8610000D";
    when 16#1760# => romdata <= X"1B3FFC00";
    when 16#1761# => romdata <= X"9A28800D";
    when 16#1762# => romdata <= X"84134001";
    when 16#1763# => romdata <= X"10BFFF3C";
    when 16#1764# => romdata <= X"C207BFFC";
    when 16#1765# => romdata <= X"C627BFE0";
    when 16#1766# => romdata <= X"A4102000";
    when 16#1767# => romdata <= X"B6102000";
    when 16#1768# => romdata <= X"AE102001";
    when 16#1769# => romdata <= X"AC103FFF";
    when 16#176A# => romdata <= X"B8102000";
    when 16#176B# => romdata <= X"C0262044";
    when 16#176C# => romdata <= X"92102000";
    when 16#176D# => romdata <= X"D127BFD4";
    when 16#176E# => romdata <= X"D327BFD0";
    when 16#176F# => romdata <= X"D527BFDC";
    when 16#1770# => romdata <= X"D727BFD8";
    when 16#1771# => romdata <= X"40000998";
    when 16#1772# => romdata <= X"90100018";
    when 16#1773# => romdata <= X"D0262040";
    when 16#1774# => romdata <= X"AA100008";
    when 16#1775# => romdata <= X"808CA0FF";
    when 16#1776# => romdata <= X"D107BFD4";
    when 16#1777# => romdata <= X"D307BFD0";
    when 16#1778# => romdata <= X"D507BFDC";
    when 16#1779# => romdata <= X"02BFFF94";
    when 16#177A# => romdata <= X"D707BFD8";
    when 16#177B# => romdata <= X"80A4E000";
    when 16#177C# => romdata <= X"0480022F";
    when 16#177D# => romdata <= X"820CE00F";
    when 16#177E# => romdata <= X"83286003";
    when 16#177F# => romdata <= X"05100032";
    when 16#1780# => romdata <= X"99A0002A";
    when 16#1781# => romdata <= X"8410A150";
    when 16#1782# => romdata <= X"9BA0002B";
    when 16#1783# => romdata <= X"D1188001";
    when 16#1784# => romdata <= X"833CE004";
    when 16#1785# => romdata <= X"80886010";
    when 16#1786# => romdata <= X"1280012A";
    when 16#1787# => romdata <= X"86102002";
    when 16#1788# => romdata <= X"80A06000";
    when 16#1789# => romdata <= X"2280000E";
    when 16#178A# => romdata <= X"91A309C8";
    when 16#178B# => romdata <= X"05100032";
    when 16#178C# => romdata <= X"8410A218";
    when 16#178D# => romdata <= X"80886001";
    when 16#178E# => romdata <= X"02800005";
    when 16#178F# => romdata <= X"83386001";
    when 16#1790# => romdata <= X"DD188000";
    when 16#1791# => romdata <= X"91A2094E";
    when 16#1792# => romdata <= X"8600E001";
    when 16#1793# => romdata <= X"80A06000";
    when 16#1794# => romdata <= X"12BFFFF9";
    when 16#1795# => romdata <= X"8400A008";
    when 16#1796# => romdata <= X"91A309C8";
    when 16#1797# => romdata <= X"C207BFF4";
    when 16#1798# => romdata <= X"80A06000";
    when 16#1799# => romdata <= X"22800020";
    when 16#179A# => romdata <= X"C627BFC4";
    when 16#179B# => romdata <= X"03100032";
    when 16#179C# => romdata <= X"D91860E0";
    when 16#179D# => romdata <= X"81AA0ACC";
    when 16#179E# => romdata <= X"01000000";
    when 16#179F# => romdata <= X"19800019";
    when 16#17A0# => romdata <= X"01000000";
    when 16#17A1# => romdata <= X"80A5A000";
    when 16#17A2# => romdata <= X"04800016";
    when 16#17A3# => romdata <= X"C407BFE0";
    when 16#17A4# => romdata <= X"80A0A000";
    when 16#17A5# => romdata <= X"048001D4";
    when 16#17A6# => romdata <= X"8600E001";
    when 16#17A7# => romdata <= X"C627BFC4";
    when 16#17A8# => romdata <= X"1B100032";
    when 16#17A9# => romdata <= X"D91B60E8";
    when 16#17AA# => romdata <= X"91A2094C";
    when 16#17AB# => romdata <= X"03100032";
    when 16#17AC# => romdata <= X"D907BFC4";
    when 16#17AD# => romdata <= X"9DA0190C";
    when 16#17AE# => romdata <= X"9DA2094E";
    when 16#17AF# => romdata <= X"D91860F0";
    when 16#17B0# => romdata <= X"A1A3884C";
    when 16#17B1# => romdata <= X"E13FBFC8";
    when 16#17B2# => romdata <= X"033F3000";
    when 16#17B3# => romdata <= X"D81FBFC8";
    when 16#17B4# => romdata <= X"9800400C";
    when 16#17B5# => romdata <= X"8204FFFF";
    when 16#17B6# => romdata <= X"10800163";
    when 16#17B7# => romdata <= X"C227BFEC";
    when 16#17B8# => romdata <= X"C627BFC4";
    when 16#17B9# => romdata <= X"03100032";
    when 16#17BA# => romdata <= X"80A5A000";
    when 16#17BB# => romdata <= X"D907BFC4";
    when 16#17BC# => romdata <= X"9DA0190C";
    when 16#17BD# => romdata <= X"9DA38948";
    when 16#17BE# => romdata <= X"D91860F0";
    when 16#17BF# => romdata <= X"A1A3884C";
    when 16#17C0# => romdata <= X"E13FBFC8";
    when 16#17C1# => romdata <= X"033F3000";
    when 16#17C2# => romdata <= X"D81FBFC8";
    when 16#17C3# => romdata <= X"12800154";
    when 16#17C4# => romdata <= X"9800400C";
    when 16#17C5# => romdata <= X"D83FBFC8";
    when 16#17C6# => romdata <= X"03100032";
    when 16#17C7# => romdata <= X"D91860F8";
    when 16#17C8# => romdata <= X"91A208CC";
    when 16#17C9# => romdata <= X"D91FBFC8";
    when 16#17CA# => romdata <= X"81AA0ACC";
    when 16#17CB# => romdata <= X"01000000";
    when 16#17CC# => romdata <= X"2D8001C3";
    when 16#17CD# => romdata <= X"C027BFEC";
    when 16#17CE# => romdata <= X"99A000AC";
    when 16#17CF# => romdata <= X"81AA0ACC";
    when 16#17D0# => romdata <= X"01000000";
    when 16#17D1# => romdata <= X"198001A8";
    when 16#17D2# => romdata <= X"01000000";
    when 16#17D3# => romdata <= X"C027BFEC";
    when 16#17D4# => romdata <= X"A2102000";
    when 16#17D5# => romdata <= X"A638001C";
    when 16#17D6# => romdata <= X"EE07BFEC";
    when 16#17D7# => romdata <= X"A4100015";
    when 16#17D8# => romdata <= X"1080010E";
    when 16#17D9# => romdata <= X"B8102000";
    when 16#17DA# => romdata <= X"80A5E000";
    when 16#17DB# => romdata <= X"1280011D";
    when 16#17DC# => romdata <= X"80A6E001";
    when 16#17DD# => romdata <= X"E207BFF0";
    when 16#17DE# => romdata <= X"F227BFE8";
    when 16#17DF# => romdata <= X"C027BFEC";
    when 16#17E0# => romdata <= X"80A6A000";
    when 16#17E1# => romdata <= X"0480000D";
    when 16#17E2# => romdata <= X"D807BFE8";
    when 16#17E3# => romdata <= X"80A32000";
    when 16#17E4# => romdata <= X"0480000A";
    when 16#17E5# => romdata <= X"80A6800C";
    when 16#17E6# => romdata <= X"04800003";
    when 16#17E7# => romdata <= X"8210001A";
    when 16#17E8# => romdata <= X"8210000C";
    when 16#17E9# => romdata <= X"DA07BFE8";
    when 16#17EA# => romdata <= X"9A234001";
    when 16#17EB# => romdata <= X"DA27BFE8";
    when 16#17EC# => romdata <= X"B4268001";
    when 16#17ED# => romdata <= X"B2264001";
    when 16#17EE# => romdata <= X"C207BFF0";
    when 16#17EF# => romdata <= X"80A06000";
    when 16#17F0# => romdata <= X"0480001B";
    when 16#17F1# => romdata <= X"80A5E000";
    when 16#17F2# => romdata <= X"0280024D";
    when 16#17F3# => romdata <= X"80A46000";
    when 16#17F4# => romdata <= X"04800013";
    when 16#17F5# => romdata <= X"D207BFEC";
    when 16#17F6# => romdata <= X"D127BFD4";
    when 16#17F7# => romdata <= X"D327BFD0";
    when 16#17F8# => romdata <= X"94100011";
    when 16#17F9# => romdata <= X"40000B0B";
    when 16#17FA# => romdata <= X"90100018";
    when 16#17FB# => romdata <= X"D027BFEC";
    when 16#17FC# => romdata <= X"94100014";
    when 16#17FD# => romdata <= X"90100018";
    when 16#17FE# => romdata <= X"40000A3B";
    when 16#17FF# => romdata <= X"D207BFEC";
    when 16#1800# => romdata <= X"92100014";
    when 16#1801# => romdata <= X"A4100008";
    when 16#1802# => romdata <= X"400007DF";
    when 16#1803# => romdata <= X"90100018";
    when 16#1804# => romdata <= X"D307BFD0";
    when 16#1805# => romdata <= X"D107BFD4";
    when 16#1806# => romdata <= X"A8100012";
    when 16#1807# => romdata <= X"C407BFF0";
    when 16#1808# => romdata <= X"94A08011";
    when 16#1809# => romdata <= X"12800252";
    when 16#180A# => romdata <= X"92100014";
    when 16#180B# => romdata <= X"D127BFD4";
    when 16#180C# => romdata <= X"D327BFD0";
    when 16#180D# => romdata <= X"90100018";
    when 16#180E# => romdata <= X"40000AB3";
    when 16#180F# => romdata <= X"92102001";
    when 16#1810# => romdata <= X"C607BFE4";
    when 16#1811# => romdata <= X"A2100008";
    when 16#1812# => romdata <= X"80A0E000";
    when 16#1813# => romdata <= X"D107BFD4";
    when 16#1814# => romdata <= X"04800009";
    when 16#1815# => romdata <= X"D307BFD0";
    when 16#1816# => romdata <= X"92100008";
    when 16#1817# => romdata <= X"94100003";
    when 16#1818# => romdata <= X"40000AEC";
    when 16#1819# => romdata <= X"90100018";
    when 16#181A# => romdata <= X"D307BFD0";
    when 16#181B# => romdata <= X"D107BFD4";
    when 16#181C# => romdata <= X"A2100008";
    when 16#181D# => romdata <= X"80A6E001";
    when 16#181E# => romdata <= X"2480013A";
    when 16#181F# => romdata <= X"D327BFC4";
    when 16#1820# => romdata <= X"C027BFF0";
    when 16#1821# => romdata <= X"DA07BFE4";
    when 16#1822# => romdata <= X"80A36000";
    when 16#1823# => romdata <= X"128001E9";
    when 16#1824# => romdata <= X"82102001";
    when 16#1825# => romdata <= X"8200401A";
    when 16#1826# => romdata <= X"8288601F";
    when 16#1827# => romdata <= X"12800170";
    when 16#1828# => romdata <= X"8410201C";
    when 16#1829# => romdata <= X"C607BFE8";
    when 16#182A# => romdata <= X"8600C002";
    when 16#182B# => romdata <= X"C627BFE8";
    when 16#182C# => romdata <= X"B4068002";
    when 16#182D# => romdata <= X"B2064002";
    when 16#182E# => romdata <= X"80A66000";
    when 16#182F# => romdata <= X"0480000A";
    when 16#1830# => romdata <= X"92100014";
    when 16#1831# => romdata <= X"D127BFD4";
    when 16#1832# => romdata <= X"D327BFD0";
    when 16#1833# => romdata <= X"94100019";
    when 16#1834# => romdata <= X"400009B8";
    when 16#1835# => romdata <= X"90100018";
    when 16#1836# => romdata <= X"D307BFD0";
    when 16#1837# => romdata <= X"D107BFD4";
    when 16#1838# => romdata <= X"A8100008";
    when 16#1839# => romdata <= X"80A6A000";
    when 16#183A# => romdata <= X"0480000A";
    when 16#183B# => romdata <= X"92100011";
    when 16#183C# => romdata <= X"D127BFD4";
    when 16#183D# => romdata <= X"D327BFD0";
    when 16#183E# => romdata <= X"9410001A";
    when 16#183F# => romdata <= X"400009AD";
    when 16#1840# => romdata <= X"90100018";
    when 16#1841# => romdata <= X"D307BFD0";
    when 16#1842# => romdata <= X"D107BFD4";
    when 16#1843# => romdata <= X"A2100008";
    when 16#1844# => romdata <= X"C807BFF4";
    when 16#1845# => romdata <= X"80A12000";
    when 16#1846# => romdata <= X"328001D3";
    when 16#1847# => romdata <= X"D127BFD4";
    when 16#1848# => romdata <= X"80A5A000";
    when 16#1849# => romdata <= X"04800200";
    when 16#184A# => romdata <= X"80A6E002";
    when 16#184B# => romdata <= X"80A5E000";
    when 16#184C# => romdata <= X"A4100015";
    when 16#184D# => romdata <= X"02800077";
    when 16#184E# => romdata <= X"AE102001";
    when 16#184F# => romdata <= X"D807BFE8";
    when 16#1850# => romdata <= X"80A32000";
    when 16#1851# => romdata <= X"0480000A";
    when 16#1852# => romdata <= X"D207BFEC";
    when 16#1853# => romdata <= X"D127BFD4";
    when 16#1854# => romdata <= X"D327BFD0";
    when 16#1855# => romdata <= X"9410000C";
    when 16#1856# => romdata <= X"40000996";
    when 16#1857# => romdata <= X"90100018";
    when 16#1858# => romdata <= X"D307BFD0";
    when 16#1859# => romdata <= X"D027BFEC";
    when 16#185A# => romdata <= X"D107BFD4";
    when 16#185B# => romdata <= X"DA07BFF0";
    when 16#185C# => romdata <= X"80A36000";
    when 16#185D# => romdata <= X"12800234";
    when 16#185E# => romdata <= X"EE07BFEC";
    when 16#185F# => romdata <= X"D327BFC4";
    when 16#1860# => romdata <= X"F807BFEC";
    when 16#1861# => romdata <= X"A4100015";
    when 16#1862# => romdata <= X"B4102001";
    when 16#1863# => romdata <= X"C607BFC4";
    when 16#1864# => romdata <= X"B208E001";
    when 16#1865# => romdata <= X"92100011";
    when 16#1866# => romdata <= X"7FFFFD24";
    when 16#1867# => romdata <= X"90100014";
    when 16#1868# => romdata <= X"90022030";
    when 16#1869# => romdata <= X"9210001C";
    when 16#186A# => romdata <= X"D027BFF4";
    when 16#186B# => romdata <= X"400007DB";
    when 16#186C# => romdata <= X"90100014";
    when 16#186D# => romdata <= X"92100011";
    when 16#186E# => romdata <= X"D027BFF0";
    when 16#186F# => romdata <= X"94100017";
    when 16#1870# => romdata <= X"4000090F";
    when 16#1871# => romdata <= X"90100018";
    when 16#1872# => romdata <= X"C402200C";
    when 16#1873# => romdata <= X"80A0A000";
    when 16#1874# => romdata <= X"82100008";
    when 16#1875# => romdata <= X"02800107";
    when 16#1876# => romdata <= X"84102001";
    when 16#1877# => romdata <= X"C427BFDC";
    when 16#1878# => romdata <= X"92100001";
    when 16#1879# => romdata <= X"40000768";
    when 16#187A# => romdata <= X"90100018";
    when 16#187B# => romdata <= X"C407BFDC";
    when 16#187C# => romdata <= X"80A0A000";
    when 16#187D# => romdata <= X"12800008";
    when 16#187E# => romdata <= X"DA07BFF0";
    when 16#187F# => romdata <= X"80A6E000";
    when 16#1880# => romdata <= X"12800006";
    when 16#1881# => romdata <= X"80A36000";
    when 16#1882# => romdata <= X"80A66000";
    when 16#1883# => romdata <= X"02800233";
    when 16#1884# => romdata <= X"C807BFF4";
    when 16#1885# => romdata <= X"80A36000";
    when 16#1886# => romdata <= X"068001E5";
    when 16#1887# => romdata <= X"80A36000";
    when 16#1888# => romdata <= X"12800008";
    when 16#1889# => romdata <= X"80A0A000";
    when 16#188A# => romdata <= X"80A6E000";
    when 16#188B# => romdata <= X"12800005";
    when 16#188C# => romdata <= X"80A0A000";
    when 16#188D# => romdata <= X"80A66000";
    when 16#188E# => romdata <= X"028001DD";
    when 16#188F# => romdata <= X"80A0A000";
    when 16#1890# => romdata <= X"1480021A";
    when 16#1891# => romdata <= X"DA07BFF4";
    when 16#1892# => romdata <= X"80A68016";
    when 16#1893# => romdata <= X"DA2C8000";
    when 16#1894# => romdata <= X"0280003C";
    when 16#1895# => romdata <= X"A404A001";
    when 16#1896# => romdata <= X"92100014";
    when 16#1897# => romdata <= X"90100018";
    when 16#1898# => romdata <= X"9410200A";
    when 16#1899# => romdata <= X"40000A31";
    when 16#189A# => romdata <= X"96102000";
    when 16#189B# => romdata <= X"80A70017";
    when 16#189C# => romdata <= X"02800106";
    when 16#189D# => romdata <= X"A8100008";
    when 16#189E# => romdata <= X"9210001C";
    when 16#189F# => romdata <= X"9410200A";
    when 16#18A0# => romdata <= X"96102000";
    when 16#18A1# => romdata <= X"40000A29";
    when 16#18A2# => romdata <= X"90100018";
    when 16#18A3# => romdata <= X"92100017";
    when 16#18A4# => romdata <= X"B8100008";
    when 16#18A5# => romdata <= X"9410200A";
    when 16#18A6# => romdata <= X"90100018";
    when 16#18A7# => romdata <= X"96102000";
    when 16#18A8# => romdata <= X"40000A22";
    when 16#18A9# => romdata <= X"B406A001";
    when 16#18AA# => romdata <= X"10BFFFBB";
    when 16#18AB# => romdata <= X"AE100008";
    when 16#18AC# => romdata <= X"B2264013";
    when 16#18AD# => romdata <= X"C627BFF0";
    when 16#18AE# => romdata <= X"10BFFE2A";
    when 16#18AF# => romdata <= X"C027BFE4";
    when 16#18B0# => romdata <= X"05100032";
    when 16#18B1# => romdata <= X"D918A238";
    when 16#18B2# => romdata <= X"99A289CC";
    when 16#18B3# => romdata <= X"8208600F";
    when 16#18B4# => romdata <= X"10BFFED4";
    when 16#18B5# => romdata <= X"86102003";
    when 16#18B6# => romdata <= X"02800152";
    when 16#18B7# => romdata <= X"88103FFF";
    when 16#18B8# => romdata <= X"A4102000";
    when 16#18B9# => romdata <= X"AE102001";
    when 16#18BA# => romdata <= X"C827BFE0";
    when 16#18BB# => romdata <= X"AC103FFF";
    when 16#18BC# => romdata <= X"10BFFEAF";
    when 16#18BD# => romdata <= X"B8102000";
    when 16#18BE# => romdata <= X"90100018";
    when 16#18BF# => romdata <= X"9410200A";
    when 16#18C0# => romdata <= X"96102000";
    when 16#18C1# => romdata <= X"40000A09";
    when 16#18C2# => romdata <= X"AE05E001";
    when 16#18C3# => romdata <= X"A8100008";
    when 16#18C4# => romdata <= X"92100011";
    when 16#18C5# => romdata <= X"7FFFFCC5";
    when 16#18C6# => romdata <= X"90100014";
    when 16#18C7# => romdata <= X"90022030";
    when 16#18C8# => romdata <= X"D027BFF4";
    when 16#18C9# => romdata <= X"80A5C016";
    when 16#18CA# => romdata <= X"D02C8000";
    when 16#18CB# => romdata <= X"92100014";
    when 16#18CC# => romdata <= X"06BFFFF2";
    when 16#18CD# => romdata <= X"A404A001";
    when 16#18CE# => romdata <= X"EE07BFEC";
    when 16#18CF# => romdata <= X"B8102000";
    when 16#18D0# => romdata <= X"92100014";
    when 16#18D1# => romdata <= X"94102001";
    when 16#18D2# => romdata <= X"4000091A";
    when 16#18D3# => romdata <= X"90100018";
    when 16#18D4# => romdata <= X"92100011";
    when 16#18D5# => romdata <= X"40000771";
    when 16#18D6# => romdata <= X"A8100008";
    when 16#18D7# => romdata <= X"80A22000";
    when 16#18D8# => romdata <= X"34800004";
    when 16#18D9# => romdata <= X"C24CBFFF";
    when 16#18DA# => romdata <= X"308001A5";
    when 16#18DB# => romdata <= X"C24CBFFF";
    when 16#18DC# => romdata <= X"80A06039";
    when 16#18DD# => romdata <= X"C40CBFFF";
    when 16#18DE# => romdata <= X"128001B0";
    when 16#18DF# => romdata <= X"8204BFFF";
    when 16#18E0# => romdata <= X"80A04015";
    when 16#18E1# => romdata <= X"32BFFFFA";
    when 16#18E2# => romdata <= X"A4100001";
    when 16#18E3# => romdata <= X"82102031";
    when 16#18E4# => romdata <= X"C22D4000";
    when 16#18E5# => romdata <= X"A604E001";
    when 16#18E6# => romdata <= X"92100011";
    when 16#18E7# => romdata <= X"400006FA";
    when 16#18E8# => romdata <= X"90100018";
    when 16#18E9# => romdata <= X"80A5E000";
    when 16#18EA# => romdata <= X"02BFFE67";
    when 16#18EB# => romdata <= X"80A70017";
    when 16#18EC# => romdata <= X"02800006";
    when 16#18ED# => romdata <= X"80A72000";
    when 16#18EE# => romdata <= X"02800004";
    when 16#18EF# => romdata <= X"9210001C";
    when 16#18F0# => romdata <= X"400006F1";
    when 16#18F1# => romdata <= X"90100018";
    when 16#18F2# => romdata <= X"92100017";
    when 16#18F3# => romdata <= X"E627BFEC";
    when 16#18F4# => romdata <= X"400006ED";
    when 16#18F5# => romdata <= X"90100018";
    when 16#18F6# => romdata <= X"10BFFD51";
    when 16#18F7# => romdata <= X"90100018";
    when 16#18F8# => romdata <= X"0480016B";
    when 16#18F9# => romdata <= X"DA07BFF0";
    when 16#18FA# => romdata <= X"8205BFFF";
    when 16#18FB# => romdata <= X"80A34001";
    when 16#18FC# => romdata <= X"16800009";
    when 16#18FD# => romdata <= X"A2234001";
    when 16#18FE# => romdata <= X"C607BFE4";
    when 16#18FF# => romdata <= X"8220400D";
    when 16#1900# => romdata <= X"84034001";
    when 16#1901# => romdata <= X"8600C001";
    when 16#1902# => romdata <= X"C427BFF0";
    when 16#1903# => romdata <= X"C627BFE4";
    when 16#1904# => romdata <= X"A2102000";
    when 16#1905# => romdata <= X"88264016";
    when 16#1906# => romdata <= X"C827BFE8";
    when 16#1907# => romdata <= X"80A5A000";
    when 16#1908# => romdata <= X"06800004";
    when 16#1909# => romdata <= X"82102000";
    when 16#190A# => romdata <= X"F227BFE8";
    when 16#190B# => romdata <= X"82100016";
    when 16#190C# => romdata <= X"D127BFD4";
    when 16#190D# => romdata <= X"D327BFD0";
    when 16#190E# => romdata <= X"B4068001";
    when 16#190F# => romdata <= X"B2064001";
    when 16#1910# => romdata <= X"90100018";
    when 16#1911# => romdata <= X"400009B0";
    when 16#1912# => romdata <= X"92102001";
    when 16#1913# => romdata <= X"D307BFD0";
    when 16#1914# => romdata <= X"D027BFEC";
    when 16#1915# => romdata <= X"10BFFECB";
    when 16#1916# => romdata <= X"D107BFD4";
    when 16#1917# => romdata <= X"E627BFEC";
    when 16#1918# => romdata <= X"84100016";
    when 16#1919# => romdata <= X"80A5E000";
    when 16#191A# => romdata <= X"228000AD";
    when 16#191B# => romdata <= X"99A01A48";
    when 16#191C# => romdata <= X"8200BFFF";
    when 16#191D# => romdata <= X"83286003";
    when 16#191E# => romdata <= X"07100032";
    when 16#191F# => romdata <= X"8610E150";
    when 16#1920# => romdata <= X"D918C001";
    when 16#1921# => romdata <= X"03100032";
    when 16#1922# => romdata <= X"DD186100";
    when 16#1923# => romdata <= X"9DA389CC";
    when 16#1924# => romdata <= X"99A01A48";
    when 16#1925# => romdata <= X"D927BFC4";
    when 16#1926# => romdata <= X"99A0190C";
    when 16#1927# => romdata <= X"99A208CC";
    when 16#1928# => romdata <= X"C607BFC4";
    when 16#1929# => romdata <= X"8200E030";
    when 16#192A# => romdata <= X"C22D4000";
    when 16#192B# => romdata <= X"D83FBFC8";
    when 16#192C# => romdata <= X"D11FBFC8";
    when 16#192D# => romdata <= X"91A388C8";
    when 16#192E# => romdata <= X"81AA0ACC";
    when 16#192F# => romdata <= X"01000000";
    when 16#1930# => romdata <= X"0DBFFD16";
    when 16#1931# => romdata <= X"A4056001";
    when 16#1932# => romdata <= X"09100032";
    when 16#1933# => romdata <= X"DD1920E0";
    when 16#1934# => romdata <= X"9DA388CC";
    when 16#1935# => romdata <= X"81AA0ACE";
    when 16#1936# => romdata <= X"01000000";
    when 16#1937# => romdata <= X"0D8000D3";
    when 16#1938# => romdata <= X"80A0A001";
    when 16#1939# => romdata <= X"04800040";
    when 16#193A# => romdata <= X"1B100032";
    when 16#193B# => romdata <= X"881120E0";
    when 16#193C# => romdata <= X"E11B60E8";
    when 16#193D# => romdata <= X"1080000A";
    when 16#193E# => romdata <= X"82102001";
    when 16#193F# => romdata <= X"DD190000";
    when 16#1940# => romdata <= X"9DA388CC";
    when 16#1941# => romdata <= X"81AB8AC8";
    when 16#1942# => romdata <= X"01000000";
    when 16#1943# => romdata <= X"29800028";
    when 16#1944# => romdata <= X"E607BFEC";
    when 16#1945# => romdata <= X"36800035";
    when 16#1946# => romdata <= X"91A0002A";
    when 16#1947# => romdata <= X"99A30950";
    when 16#1948# => romdata <= X"9DA01A4C";
    when 16#1949# => romdata <= X"DD27BFC4";
    when 16#194A# => romdata <= X"9DA0190E";
    when 16#194B# => romdata <= X"99A308CE";
    when 16#194C# => romdata <= X"91A20950";
    when 16#194D# => romdata <= X"82006001";
    when 16#194E# => romdata <= X"81AB0AC8";
    when 16#194F# => romdata <= X"80A04002";
    when 16#1950# => romdata <= X"D807BFC4";
    when 16#1951# => romdata <= X"86032030";
    when 16#1952# => romdata <= X"C62C8000";
    when 16#1953# => romdata <= X"01000000";
    when 16#1954# => romdata <= X"19BFFFEB";
    when 16#1955# => romdata <= X"A404A001";
    when 16#1956# => romdata <= X"10BFFCF1";
    when 16#1957# => romdata <= X"90100018";
    when 16#1958# => romdata <= X"C807BFC4";
    when 16#1959# => romdata <= X"80A12000";
    when 16#195A# => romdata <= X"32BFFEC7";
    when 16#195B# => romdata <= X"C027BFF0";
    when 16#195C# => romdata <= X"D127BFC4";
    when 16#195D# => romdata <= X"053FFC00";
    when 16#195E# => romdata <= X"C207BFC4";
    when 16#195F# => romdata <= X"80A84002";
    when 16#1960# => romdata <= X"32BFFEC1";
    when 16#1961# => romdata <= X"C027BFF0";
    when 16#1962# => romdata <= X"051FFC00";
    when 16#1963# => romdata <= X"80884002";
    when 16#1964# => romdata <= X"22BFFEBD";
    when 16#1965# => romdata <= X"C027BFF0";
    when 16#1966# => romdata <= X"98102001";
    when 16#1967# => romdata <= X"B2066001";
    when 16#1968# => romdata <= X"B406A001";
    when 16#1969# => romdata <= X"10BFFEB8";
    when 16#196A# => romdata <= X"D827BFF0";
    when 16#196B# => romdata <= X"C24CBFFF";
    when 16#196C# => romdata <= X"80A06039";
    when 16#196D# => romdata <= X"C40CBFFF";
    when 16#196E# => romdata <= X"12BFFCD5";
    when 16#196F# => romdata <= X"8204BFFF";
    when 16#1970# => romdata <= X"80A04015";
    when 16#1971# => romdata <= X"32BFFFFA";
    when 16#1972# => romdata <= X"A4100001";
    when 16#1973# => romdata <= X"82102030";
    when 16#1974# => romdata <= X"A604E001";
    when 16#1975# => romdata <= X"C22D4000";
    when 16#1976# => romdata <= X"84102031";
    when 16#1977# => romdata <= X"10BFFCCD";
    when 16#1978# => romdata <= X"82100015";
    when 16#1979# => romdata <= X"91A0002A";
    when 16#197A# => romdata <= X"10BFFD93";
    when 16#197B# => romdata <= X"93A0002B";
    when 16#197C# => romdata <= X"92100001";
    when 16#197D# => romdata <= X"C227BFDC";
    when 16#197E# => romdata <= X"400006C8";
    when 16#197F# => romdata <= X"90100014";
    when 16#1980# => romdata <= X"C207BFDC";
    when 16#1981# => romdata <= X"10BFFEF6";
    when 16#1982# => romdata <= X"84100008";
    when 16#1983# => romdata <= X"80A72000";
    when 16#1984# => romdata <= X"36BFFD95";
    when 16#1985# => romdata <= X"95A209CC";
    when 16#1986# => romdata <= X"80A5A000";
    when 16#1987# => romdata <= X"12BFFE4C";
    when 16#1988# => romdata <= X"03100032";
    when 16#1989# => romdata <= X"D51860F8";
    when 16#198A# => romdata <= X"99A3094A";
    when 16#198B# => romdata <= X"81AB0AC8";
    when 16#198C# => romdata <= X"01000000";
    when 16#198D# => romdata <= X"17BFFE47";
    when 16#198E# => romdata <= X"C027BFEC";
    when 16#198F# => romdata <= X"A2102000";
    when 16#1990# => romdata <= X"EE07BFEC";
    when 16#1991# => romdata <= X"82102031";
    when 16#1992# => romdata <= X"A604E001";
    when 16#1993# => romdata <= X"C22D4000";
    when 16#1994# => romdata <= X"A4056001";
    when 16#1995# => romdata <= X"10BFFF51";
    when 16#1996# => romdata <= X"B8102000";
    when 16#1997# => romdata <= X"84102020";
    when 16#1998# => romdata <= X"82208001";
    when 16#1999# => romdata <= X"80A06004";
    when 16#199A# => romdata <= X"04800133";
    when 16#199B# => romdata <= X"C407BFE8";
    when 16#199C# => romdata <= X"82007FFC";
    when 16#199D# => romdata <= X"84008001";
    when 16#199E# => romdata <= X"B4068001";
    when 16#199F# => romdata <= X"B2064001";
    when 16#19A0# => romdata <= X"10BFFE8E";
    when 16#19A1# => romdata <= X"C427BFE8";
    when 16#19A2# => romdata <= X"9210001C";
    when 16#19A3# => romdata <= X"90100018";
    when 16#19A4# => romdata <= X"9410200A";
    when 16#19A5# => romdata <= X"96102000";
    when 16#19A6# => romdata <= X"40000924";
    when 16#19A7# => romdata <= X"B406A001";
    when 16#19A8# => romdata <= X"B8100008";
    when 16#19A9# => romdata <= X"10BFFEBC";
    when 16#19AA# => romdata <= X"AE100008";
    when 16#19AB# => romdata <= X"91A0002A";
    when 16#19AC# => romdata <= X"93A0002B";
    when 16#19AD# => romdata <= X"82A00013";
    when 16#19AE# => romdata <= X"02BFFDE9";
    when 16#19AF# => romdata <= X"86102002";
    when 16#19B0# => romdata <= X"8408600F";
    when 16#19B1# => romdata <= X"07100032";
    when 16#19B2# => romdata <= X"8528A003";
    when 16#19B3# => romdata <= X"8610E150";
    when 16#19B4# => romdata <= X"D118C002";
    when 16#19B5# => romdata <= X"83386004";
    when 16#19B6# => romdata <= X"91A28948";
    when 16#19B7# => romdata <= X"80A06000";
    when 16#19B8# => romdata <= X"02BFFDDF";
    when 16#19B9# => romdata <= X"86102002";
    when 16#19BA# => romdata <= X"05100032";
    when 16#19BB# => romdata <= X"8410A218";
    when 16#19BC# => romdata <= X"80886001";
    when 16#19BD# => romdata <= X"02800005";
    when 16#19BE# => romdata <= X"83386001";
    when 16#19BF# => romdata <= X"D9188000";
    when 16#19C0# => romdata <= X"91A2094C";
    when 16#19C1# => romdata <= X"8600E001";
    when 16#19C2# => romdata <= X"80A06000";
    when 16#19C3# => romdata <= X"12BFFFF9";
    when 16#19C4# => romdata <= X"8400A008";
    when 16#19C5# => romdata <= X"10BFFDD3";
    when 16#19C6# => romdata <= X"C207BFF4";
    when 16#19C7# => romdata <= X"D927BFC4";
    when 16#19C8# => romdata <= X"99A0190C";
    when 16#19C9# => romdata <= X"91A208CC";
    when 16#19CA# => romdata <= X"80A0A001";
    when 16#19CB# => romdata <= X"A4056001";
    when 16#19CC# => romdata <= X"C607BFC4";
    when 16#19CD# => romdata <= X"8200E030";
    when 16#19CE# => romdata <= X"07100032";
    when 16#19CF# => romdata <= X"8610E150";
    when 16#19D0# => romdata <= X"C22D4000";
    when 16#19D1# => romdata <= X"D83FBFC8";
    when 16#19D2# => romdata <= X"8200BFFF";
    when 16#19D3# => romdata <= X"83286003";
    when 16#19D4# => romdata <= X"E118C001";
    when 16#19D5# => romdata <= X"DD1FBFC8";
    when 16#19D6# => romdata <= X"02800012";
    when 16#19D7# => romdata <= X"A1A4094E";
    when 16#19D8# => romdata <= X"1B100032";
    when 16#19D9# => romdata <= X"DD1B60E8";
    when 16#19DA# => romdata <= X"82102001";
    when 16#19DB# => romdata <= X"91A2094E";
    when 16#19DC# => romdata <= X"99A01A48";
    when 16#19DD# => romdata <= X"D927BFC4";
    when 16#19DE# => romdata <= X"99A0190C";
    when 16#19DF# => romdata <= X"C807BFC4";
    when 16#19E0# => romdata <= X"86012030";
    when 16#19E1# => romdata <= X"C62D4001";
    when 16#19E2# => romdata <= X"82006001";
    when 16#19E3# => romdata <= X"80A04002";
    when 16#19E4# => romdata <= X"12BFFFF7";
    when 16#19E5# => romdata <= X"91A208CC";
    when 16#19E6# => romdata <= X"82007FFF";
    when 16#19E7# => romdata <= X"A4048001";
    when 16#19E8# => romdata <= X"03100032";
    when 16#19E9# => romdata <= X"D9186100";
    when 16#19EA# => romdata <= X"9DA4084C";
    when 16#19EB# => romdata <= X"81AA0ACE";
    when 16#19EC# => romdata <= X"01000000";
    when 16#19ED# => romdata <= X"2DBFFF7E";
    when 16#19EE# => romdata <= X"E607BFEC";
    when 16#19EF# => romdata <= X"99A308D0";
    when 16#19F0# => romdata <= X"81AA0ACC";
    when 16#19F1# => romdata <= X"01000000";
    when 16#19F2# => romdata <= X"19BFFF87";
    when 16#19F3# => romdata <= X"01000000";
    when 16#19F4# => romdata <= X"10800004";
    when 16#19F5# => romdata <= X"C24CBFFF";
    when 16#19F6# => romdata <= X"A4100001";
    when 16#19F7# => romdata <= X"C24CBFFF";
    when 16#19F8# => romdata <= X"80A06030";
    when 16#19F9# => romdata <= X"02BFFFFD";
    when 16#19FA# => romdata <= X"8204BFFF";
    when 16#19FB# => romdata <= X"10BFFC4C";
    when 16#19FC# => romdata <= X"90100018";
    when 16#19FD# => romdata <= X"05100032";
    when 16#19FE# => romdata <= X"DD18A0B8";
    when 16#19FF# => romdata <= X"10BFFC97";
    when 16#1A00# => romdata <= X"99A3084E";
    when 16#1A01# => romdata <= X"AE102001";
    when 16#1A02# => romdata <= X"80A72000";
    when 16#1A03# => romdata <= X"04800037";
    when 16#1A04# => romdata <= X"8810001C";
    when 16#1A05# => romdata <= X"F827BFE0";
    when 16#1A06# => romdata <= X"10BFFCEA";
    when 16#1A07# => romdata <= X"AC10001C";
    when 16#1A08# => romdata <= X"10BFFFFA";
    when 16#1A09# => romdata <= X"AE102000";
    when 16#1A0A# => romdata <= X"10BFFF61";
    when 16#1A0B# => romdata <= X"E607BFEC";
    when 16#1A0C# => romdata <= X"C2046010";
    when 16#1A0D# => romdata <= X"82006003";
    when 16#1A0E# => romdata <= X"83286002";
    when 16#1A0F# => romdata <= X"82044001";
    when 16#1A10# => romdata <= X"D0006004";
    when 16#1A11# => romdata <= X"D127BFD4";
    when 16#1A12# => romdata <= X"400005DA";
    when 16#1A13# => romdata <= X"D327BFD0";
    when 16#1A14# => romdata <= X"82102020";
    when 16#1A15# => romdata <= X"D307BFD0";
    when 16#1A16# => romdata <= X"82204008";
    when 16#1A17# => romdata <= X"10BFFE0E";
    when 16#1A18# => romdata <= X"D107BFD4";
    when 16#1A19# => romdata <= X"D327BFD0";
    when 16#1A1A# => romdata <= X"90100014";
    when 16#1A1B# => romdata <= X"4000062B";
    when 16#1A1C# => romdata <= X"92100011";
    when 16#1A1D# => romdata <= X"D107BFD4";
    when 16#1A1E# => romdata <= X"80A22000";
    when 16#1A1F# => romdata <= X"16BFFE29";
    when 16#1A20# => romdata <= X"D307BFD0";
    when 16#1A21# => romdata <= X"92100014";
    when 16#1A22# => romdata <= X"90100018";
    when 16#1A23# => romdata <= X"9410200A";
    when 16#1A24# => romdata <= X"400008A6";
    when 16#1A25# => romdata <= X"96102000";
    when 16#1A26# => romdata <= X"A604FFFF";
    when 16#1A27# => romdata <= X"A8100008";
    when 16#1A28# => romdata <= X"80A5E000";
    when 16#1A29# => romdata <= X"EC07BFE0";
    when 16#1A2A# => romdata <= X"D107BFD4";
    when 16#1A2B# => romdata <= X"02BFFE1D";
    when 16#1A2C# => romdata <= X"D307BFD0";
    when 16#1A2D# => romdata <= X"D207BFEC";
    when 16#1A2E# => romdata <= X"90100018";
    when 16#1A2F# => romdata <= X"9410200A";
    when 16#1A30# => romdata <= X"4000089A";
    when 16#1A31# => romdata <= X"96102000";
    when 16#1A32# => romdata <= X"D307BFD0";
    when 16#1A33# => romdata <= X"D027BFEC";
    when 16#1A34# => romdata <= X"10BFFE14";
    when 16#1A35# => romdata <= X"D107BFD4";
    when 16#1A36# => romdata <= X"80A5A00F";
    when 16#1A37# => romdata <= X"82402000";
    when 16#1A38# => romdata <= X"10BFFD33";
    when 16#1A39# => romdata <= X"A40C8001";
    when 16#1A3A# => romdata <= X"98102001";
    when 16#1A3B# => romdata <= X"AC102001";
    when 16#1A3C# => romdata <= X"D827BFE0";
    when 16#1A3D# => romdata <= X"10BFFD2E";
    when 16#1A3E# => romdata <= X"B8102001";
    when 16#1A3F# => romdata <= X"D407BFF0";
    when 16#1A40# => romdata <= X"92100014";
    when 16#1A41# => romdata <= X"D127BFD4";
    when 16#1A42# => romdata <= X"D327BFD0";
    when 16#1A43# => romdata <= X"400008C1";
    when 16#1A44# => romdata <= X"90100018";
    when 16#1A45# => romdata <= X"D307BFD0";
    when 16#1A46# => romdata <= X"A8100008";
    when 16#1A47# => romdata <= X"10BFFDC4";
    when 16#1A48# => romdata <= X"D107BFD4";
    when 16#1A49# => romdata <= X"04BFFE03";
    when 16#1A4A# => romdata <= X"80A5E000";
    when 16#1A4B# => romdata <= X"80A5A000";
    when 16#1A4C# => romdata <= X"12BFFD89";
    when 16#1A4D# => romdata <= X"92100011";
    when 16#1A4E# => romdata <= X"94102005";
    when 16#1A4F# => romdata <= X"96102000";
    when 16#1A50# => romdata <= X"4000087A";
    when 16#1A51# => romdata <= X"90100018";
    when 16#1A52# => romdata <= X"A2100008";
    when 16#1A53# => romdata <= X"90100014";
    when 16#1A54# => romdata <= X"400005F2";
    when 16#1A55# => romdata <= X"92100011";
    when 16#1A56# => romdata <= X"80A22000";
    when 16#1A57# => romdata <= X"34BFFF3A";
    when 16#1A58# => romdata <= X"EE07BFEC";
    when 16#1A59# => romdata <= X"10BFFD7D";
    when 16#1A5A# => romdata <= X"A638001C";
    when 16#1A5B# => romdata <= X"D127BFD4";
    when 16#1A5C# => romdata <= X"D327BFD0";
    when 16#1A5D# => romdata <= X"400008A7";
    when 16#1A5E# => romdata <= X"90100018";
    when 16#1A5F# => romdata <= X"D107BFD4";
    when 16#1A60# => romdata <= X"A8100008";
    when 16#1A61# => romdata <= X"10BFFDAA";
    when 16#1A62# => romdata <= X"D307BFD0";
    when 16#1A63# => romdata <= X"D807BFE8";
    when 16#1A64# => romdata <= X"80A32000";
    when 16#1A65# => romdata <= X"22800040";
    when 16#1A66# => romdata <= X"C207BFFC";
    when 16#1A67# => romdata <= X"82006433";
    when 16#1A68# => romdata <= X"E207BFF0";
    when 16#1A69# => romdata <= X"10BFFEA3";
    when 16#1A6A# => romdata <= X"F227BFE8";
    when 16#1A6B# => romdata <= X"80A0A000";
    when 16#1A6C# => romdata <= X"0480000F";
    when 16#1A6D# => romdata <= X"92100014";
    when 16#1A6E# => romdata <= X"94102001";
    when 16#1A6F# => romdata <= X"4000077D";
    when 16#1A70# => romdata <= X"90100018";
    when 16#1A71# => romdata <= X"92100011";
    when 16#1A72# => romdata <= X"400005D4";
    when 16#1A73# => romdata <= X"A8100008";
    when 16#1A74# => romdata <= X"80A22000";
    when 16#1A75# => romdata <= X"0480004B";
    when 16#1A76# => romdata <= X"C407BFF4";
    when 16#1A77# => romdata <= X"80A0A039";
    when 16#1A78# => romdata <= X"0280003A";
    when 16#1A79# => romdata <= X"8400A001";
    when 16#1A7A# => romdata <= X"C427BFF4";
    when 16#1A7B# => romdata <= X"C607BFF4";
    when 16#1A7C# => romdata <= X"C62C8000";
    when 16#1A7D# => romdata <= X"10BFFE69";
    when 16#1A7E# => romdata <= X"A404A001";
    when 16#1A7F# => romdata <= X"3280000A";
    when 16#1A80# => romdata <= X"C24CBFFF";
    when 16#1A81# => romdata <= X"C207BFF4";
    when 16#1A82# => romdata <= X"80886001";
    when 16#1A83# => romdata <= X"12BFFE59";
    when 16#1A84# => romdata <= X"C24CBFFF";
    when 16#1A85# => romdata <= X"10800005";
    when 16#1A86# => romdata <= X"80A06030";
    when 16#1A87# => romdata <= X"A4100001";
    when 16#1A88# => romdata <= X"C24CBFFF";
    when 16#1A89# => romdata <= X"80A06030";
    when 16#1A8A# => romdata <= X"02BFFFFD";
    when 16#1A8B# => romdata <= X"8204BFFF";
    when 16#1A8C# => romdata <= X"10BFFE5B";
    when 16#1A8D# => romdata <= X"92100011";
    when 16#1A8E# => romdata <= X"8400A001";
    when 16#1A8F# => romdata <= X"10BFFE57";
    when 16#1A90# => romdata <= X"C4284000";
    when 16#1A91# => romdata <= X"D205E004";
    when 16#1A92# => romdata <= X"D327BFD0";
    when 16#1A93# => romdata <= X"D127BFD4";
    when 16#1A94# => romdata <= X"40000675";
    when 16#1A95# => romdata <= X"90100018";
    when 16#1A96# => romdata <= X"C407BFEC";
    when 16#1A97# => romdata <= X"D400A010";
    when 16#1A98# => romdata <= X"9200A00C";
    when 16#1A99# => romdata <= X"A4100008";
    when 16#1A9A# => romdata <= X"9402A002";
    when 16#1A9B# => romdata <= X"9002200C";
    when 16#1A9C# => romdata <= X"4000047B";
    when 16#1A9D# => romdata <= X"952AA002";
    when 16#1A9E# => romdata <= X"90100018";
    when 16#1A9F# => romdata <= X"92100012";
    when 16#1AA0# => romdata <= X"4000074C";
    when 16#1AA1# => romdata <= X"94102001";
    when 16#1AA2# => romdata <= X"D307BFD0";
    when 16#1AA3# => romdata <= X"10BFFDBC";
    when 16#1AA4# => romdata <= X"AE100008";
    when 16#1AA5# => romdata <= X"84102036";
    when 16#1AA6# => romdata <= X"E207BFF0";
    when 16#1AA7# => romdata <= X"82208001";
    when 16#1AA8# => romdata <= X"10BFFE64";
    when 16#1AA9# => romdata <= X"F227BFE8";
    when 16#1AAA# => romdata <= X"C807BFF4";
    when 16#1AAB# => romdata <= X"80A12039";
    when 16#1AAC# => romdata <= X"02800006";
    when 16#1AAD# => romdata <= X"D807BFF4";
    when 16#1AAE# => romdata <= X"82032001";
    when 16#1AAF# => romdata <= X"C22C8000";
    when 16#1AB0# => romdata <= X"10BFFE36";
    when 16#1AB1# => romdata <= X"A404A001";
    when 16#1AB2# => romdata <= X"82102039";
    when 16#1AB3# => romdata <= X"C22C8000";
    when 16#1AB4# => romdata <= X"10BFFE27";
    when 16#1AB5# => romdata <= X"A404A001";
    when 16#1AB6# => romdata <= X"80A12039";
    when 16#1AB7# => romdata <= X"02BFFFFB";
    when 16#1AB8# => romdata <= X"D807BFF0";
    when 16#1AB9# => romdata <= X"833B201F";
    when 16#1ABA# => romdata <= X"8220400C";
    when 16#1ABB# => romdata <= X"8330601F";
    when 16#1ABC# => romdata <= X"88010001";
    when 16#1ABD# => romdata <= X"C82C8000";
    when 16#1ABE# => romdata <= X"10BFFE28";
    when 16#1ABF# => romdata <= X"A404A001";
    when 16#1AC0# => romdata <= X"12BFFFBC";
    when 16#1AC1# => romdata <= X"C607BFF4";
    when 16#1AC2# => romdata <= X"C207BFF4";
    when 16#1AC3# => romdata <= X"80886001";
    when 16#1AC4# => romdata <= X"22BFFFB9";
    when 16#1AC5# => romdata <= X"C62C8000";
    when 16#1AC6# => romdata <= X"10BFFFB1";
    when 16#1AC7# => romdata <= X"C407BFF4";
    when 16#1AC8# => romdata <= X"80A5A00F";
    when 16#1AC9# => romdata <= X"92102000";
    when 16#1ACA# => romdata <= X"82402000";
    when 16#1ACB# => romdata <= X"10BFFCA2";
    when 16#1ACC# => romdata <= X"A4084012";
    when 16#1ACD# => romdata <= X"02BFFD62";
    when 16#1ACE# => romdata <= X"80A66000";
    when 16#1ACF# => romdata <= X"10BFFD5A";
    when 16#1AD0# => romdata <= X"8400601C";
    when 16#1AD1# => romdata <= X"9DE3BFA0";
    when 16#1AD2# => romdata <= X"80A62000";
    when 16#1AD3# => romdata <= X"02800050";
    when 16#1AD4# => romdata <= X"03100031";
    when 16#1AD5# => romdata <= X"C216200C";
    when 16#1AD6# => romdata <= X"80886200";
    when 16#1AD7# => romdata <= X"02800044";
    when 16#1AD8# => romdata <= X"01000000";
    when 16#1AD9# => romdata <= X"03100032";
    when 16#1ADA# => romdata <= X"D00062C8";
    when 16#1ADB# => romdata <= X"80A22000";
    when 16#1ADC# => romdata <= X"22800007";
    when 16#1ADD# => romdata <= X"C616200C";
    when 16#1ADE# => romdata <= X"C2022038";
    when 16#1ADF# => romdata <= X"80A06000";
    when 16#1AE0# => romdata <= X"0280003F";
    when 16#1AE1# => romdata <= X"01000000";
    when 16#1AE2# => romdata <= X"C616200C";
    when 16#1AE3# => romdata <= X"8328E010";
    when 16#1AE4# => romdata <= X"85386010";
    when 16#1AE5# => romdata <= X"8088A008";
    when 16#1AE6# => romdata <= X"22800028";
    when 16#1AE7# => romdata <= X"83306010";
    when 16#1AE8# => romdata <= X"E2062010";
    when 16#1AE9# => romdata <= X"80A46000";
    when 16#1AEA# => romdata <= X"02800023";
    when 16#1AEB# => romdata <= X"8088A003";
    when 16#1AEC# => romdata <= X"E0060000";
    when 16#1AED# => romdata <= X"E2260000";
    when 16#1AEE# => romdata <= X"A0240011";
    when 16#1AEF# => romdata <= X"12800003";
    when 16#1AF0# => romdata <= X"82102000";
    when 16#1AF1# => romdata <= X"C2062014";
    when 16#1AF2# => romdata <= X"80A42000";
    when 16#1AF3# => romdata <= X"14800008";
    when 16#1AF4# => romdata <= X"C2262008";
    when 16#1AF5# => romdata <= X"1080001F";
    when 16#1AF6# => romdata <= X"8088E200";
    when 16#1AF7# => romdata <= X"A0240008";
    when 16#1AF8# => romdata <= X"80A42000";
    when 16#1AF9# => romdata <= X"2480001A";
    when 16#1AFA# => romdata <= X"C616200C";
    when 16#1AFB# => romdata <= X"C2062024";
    when 16#1AFC# => romdata <= X"D006201C";
    when 16#1AFD# => romdata <= X"92100011";
    when 16#1AFE# => romdata <= X"9FC04000";
    when 16#1AFF# => romdata <= X"94100010";
    when 16#1B00# => romdata <= X"80A22000";
    when 16#1B01# => romdata <= X"14BFFFF6";
    when 16#1B02# => romdata <= X"A2044008";
    when 16#1B03# => romdata <= X"C416200C";
    when 16#1B04# => romdata <= X"8410A040";
    when 16#1B05# => romdata <= X"82103FFF";
    when 16#1B06# => romdata <= X"8088A200";
    when 16#1B07# => romdata <= X"1280000A";
    when 16#1B08# => romdata <= X"C436200C";
    when 16#1B09# => romdata <= X"40000FB1";
    when 16#1B0A# => romdata <= X"90062058";
    when 16#1B0B# => romdata <= X"10800006";
    when 16#1B0C# => romdata <= X"82103FFF";
    when 16#1B0D# => romdata <= X"83306010";
    when 16#1B0E# => romdata <= X"80886200";
    when 16#1B0F# => romdata <= X"02800007";
    when 16#1B10# => romdata <= X"82102000";
    when 16#1B11# => romdata <= X"81C7E008";
    when 16#1B12# => romdata <= X"91E80001";
    when 16#1B13# => romdata <= X"8088E200";
    when 16#1B14# => romdata <= X"12BFFFFD";
    when 16#1B15# => romdata <= X"82102000";
    when 16#1B16# => romdata <= X"40000FA4";
    when 16#1B17# => romdata <= X"90062058";
    when 16#1B18# => romdata <= X"82102000";
    when 16#1B19# => romdata <= X"81C7E008";
    when 16#1B1A# => romdata <= X"91E80001";
    when 16#1B1B# => romdata <= X"40000F89";
    when 16#1B1C# => romdata <= X"90062058";
    when 16#1B1D# => romdata <= X"10BFFFBD";
    when 16#1B1E# => romdata <= X"03100032";
    when 16#1B1F# => romdata <= X"40000067";
    when 16#1B20# => romdata <= X"01000000";
    when 16#1B21# => romdata <= X"10BFFFC2";
    when 16#1B22# => romdata <= X"C616200C";
    when 16#1B23# => romdata <= X"F00063FC";
    when 16#1B24# => romdata <= X"0310001A";
    when 16#1B25# => romdata <= X"400002FA";
    when 16#1B26# => romdata <= X"93E86344";
    when 16#1B27# => romdata <= X"01000000";
    when 16#1B28# => romdata <= X"13100026";
    when 16#1B29# => romdata <= X"92126148";
    when 16#1B2A# => romdata <= X"8213C000";
    when 16#1B2B# => romdata <= X"400002F4";
    when 16#1B2C# => romdata <= X"9E104000";
    when 16#1B2D# => romdata <= X"01000000";
    when 16#1B2E# => romdata <= X"03100031";
    when 16#1B2F# => romdata <= X"D00063FC";
    when 16#1B30# => romdata <= X"8213C000";
    when 16#1B31# => romdata <= X"7FFFFFF7";
    when 16#1B32# => romdata <= X"9E104000";
    when 16#1B33# => romdata <= X"01000000";
    when 16#1B34# => romdata <= X"9DE3BFA0";
    when 16#1B35# => romdata <= X"C216200C";
    when 16#1B36# => romdata <= X"80886200";
    when 16#1B37# => romdata <= X"12800004";
    when 16#1B38# => romdata <= X"01000000";
    when 16#1B39# => romdata <= X"40000F81";
    when 16#1B3A# => romdata <= X"90062058";
    when 16#1B3B# => romdata <= X"81C7E008";
    when 16#1B3C# => romdata <= X"91E82000";
    when 16#1B3D# => romdata <= X"11100035";
    when 16#1B3E# => romdata <= X"901220A4";
    when 16#1B3F# => romdata <= X"8213C000";
    when 16#1B40# => romdata <= X"40000F7A";
    when 16#1B41# => romdata <= X"9E104000";
    when 16#1B42# => romdata <= X"01000000";
    when 16#1B43# => romdata <= X"9DE3BFA0";
    when 16#1B44# => romdata <= X"03100032";
    when 16#1B45# => romdata <= X"D00062C8";
    when 16#1B46# => romdata <= X"1310001B";
    when 16#1B47# => romdata <= X"400002D8";
    when 16#1B48# => romdata <= X"921260D0";
    when 16#1B49# => romdata <= X"7FFFFFF4";
    when 16#1B4A# => romdata <= X"81E80000";
    when 16#1B4B# => romdata <= X"01000000";
    when 16#1B4C# => romdata <= X"9DE3BFA0";
    when 16#1B4D# => romdata <= X"C216200C";
    when 16#1B4E# => romdata <= X"80886200";
    when 16#1B4F# => romdata <= X"12800004";
    when 16#1B50# => romdata <= X"01000000";
    when 16#1B51# => romdata <= X"40000F53";
    when 16#1B52# => romdata <= X"90062058";
    when 16#1B53# => romdata <= X"81C7E008";
    when 16#1B54# => romdata <= X"91E82000";
    when 16#1B55# => romdata <= X"11100035";
    when 16#1B56# => romdata <= X"901220A4";
    when 16#1B57# => romdata <= X"8213C000";
    when 16#1B58# => romdata <= X"40000F4C";
    when 16#1B59# => romdata <= X"9E104000";
    when 16#1B5A# => romdata <= X"01000000";
    when 16#1B5B# => romdata <= X"9DE3BFA0";
    when 16#1B5C# => romdata <= X"7FFFFFF9";
    when 16#1B5D# => romdata <= X"3310001B";
    when 16#1B5E# => romdata <= X"03100032";
    when 16#1B5F# => romdata <= X"F00062C8";
    when 16#1B60# => romdata <= X"400002BF";
    when 16#1B61# => romdata <= X"93EE6130";
    when 16#1B62# => romdata <= X"01000000";
    when 16#1B63# => romdata <= X"9DE3BF90";
    when 16#1B64# => romdata <= X"03100025";
    when 16#1B65# => romdata <= X"821061CC";
    when 16#1B66# => romdata <= X"C2262020";
    when 16#1B67# => romdata <= X"03100025";
    when 16#1B68# => romdata <= X"82106174";
    when 16#1B69# => romdata <= X"C2262024";
    when 16#1B6A# => romdata <= X"03100025";
    when 16#1B6B# => romdata <= X"8210611C";
    when 16#1B6C# => romdata <= X"F026201C";
    when 16#1B6D# => romdata <= X"C2262028";
    when 16#1B6E# => romdata <= X"F236200C";
    when 16#1B6F# => romdata <= X"F436200E";
    when 16#1B70# => romdata <= X"C0260000";
    when 16#1B71# => romdata <= X"C0262004";
    when 16#1B72# => romdata <= X"C0262008";
    when 16#1B73# => romdata <= X"C0262010";
    when 16#1B74# => romdata <= X"C0262014";
    when 16#1B75# => romdata <= X"C0262018";
    when 16#1B76# => romdata <= X"03100025";
    when 16#1B77# => romdata <= X"82106100";
    when 16#1B78# => romdata <= X"C226202C";
    when 16#1B79# => romdata <= X"A007BFF4";
    when 16#1B7A# => romdata <= X"40000F4B";
    when 16#1B7B# => romdata <= X"90100010";
    when 16#1B7C# => romdata <= X"90100010";
    when 16#1B7D# => romdata <= X"40000F5E";
    when 16#1B7E# => romdata <= X"92102001";
    when 16#1B7F# => romdata <= X"92100010";
    when 16#1B80# => romdata <= X"40000F0C";
    when 16#1B81# => romdata <= X"90062058";
    when 16#1B82# => romdata <= X"40000F4E";
    when 16#1B83# => romdata <= X"90100010";
    when 16#1B84# => romdata <= X"81C7E008";
    when 16#1B85# => romdata <= X"81E80000";
    when 16#1B86# => romdata <= X"9DE3BFA0";
    when 16#1B87# => romdata <= X"0310001B";
    when 16#1B88# => romdata <= X"821060A0";
    when 16#1B89# => romdata <= X"C226203C";
    when 16#1B8A# => romdata <= X"82102001";
    when 16#1B8B# => romdata <= X"C2262038";
    when 16#1B8C# => romdata <= X"82102003";
    when 16#1B8D# => romdata <= X"D0062004";
    when 16#1B8E# => romdata <= X"C22622E4";
    when 16#1B8F# => romdata <= X"C02622E0";
    when 16#1B90# => romdata <= X"820622EC";
    when 16#1B91# => romdata <= X"C22622E8";
    when 16#1B92# => romdata <= X"96100018";
    when 16#1B93# => romdata <= X"92102006";
    when 16#1B94# => romdata <= X"7FFFFFCF";
    when 16#1B95# => romdata <= X"94102000";
    when 16#1B96# => romdata <= X"D0062008";
    when 16#1B97# => romdata <= X"96100018";
    when 16#1B98# => romdata <= X"B6100018";
    when 16#1B99# => romdata <= X"9210200A";
    when 16#1B9A# => romdata <= X"7FFFFFC9";
    when 16#1B9B# => romdata <= X"94102001";
    when 16#1B9C# => romdata <= X"F006200C";
    when 16#1B9D# => romdata <= X"B210200A";
    when 16#1B9E# => romdata <= X"7FFFFFC5";
    when 16#1B9F# => romdata <= X"95E82002";
    when 16#1BA0# => romdata <= X"01000000";
    when 16#1BA1# => romdata <= X"9DE3BFA0";
    when 16#1BA2# => romdata <= X"832E6002";
    when 16#1BA3# => romdata <= X"A12E6004";
    when 16#1BA4# => romdata <= X"A0240001";
    when 16#1BA5# => romdata <= X"832C2004";
    when 16#1BA6# => romdata <= X"90100018";
    when 16#1BA7# => romdata <= X"A0040001";
    when 16#1BA8# => romdata <= X"7FFFEE81";
    when 16#1BA9# => romdata <= X"9204200C";
    when 16#1BAA# => romdata <= X"B0922000";
    when 16#1BAB# => romdata <= X"02800008";
    when 16#1BAC# => romdata <= X"9006200C";
    when 16#1BAD# => romdata <= X"F2262004";
    when 16#1BAE# => romdata <= X"C0260000";
    when 16#1BAF# => romdata <= X"D0262008";
    when 16#1BB0# => romdata <= X"94100010";
    when 16#1BB1# => romdata <= X"400003F9";
    when 16#1BB2# => romdata <= X"92102000";
    when 16#1BB3# => romdata <= X"81C7E008";
    when 16#1BB4# => romdata <= X"81E80000";
    when 16#1BB5# => romdata <= X"9DE3BF90";
    when 16#1BB6# => romdata <= X"7FFFFF9F";
    when 16#1BB7# => romdata <= X"01000000";
    when 16#1BB8# => romdata <= X"03100031";
    when 16#1BB9# => romdata <= X"E20063FC";
    when 16#1BBA# => romdata <= X"C2046038";
    when 16#1BBB# => romdata <= X"80A06000";
    when 16#1BBC# => romdata <= X"02800032";
    when 16#1BBD# => romdata <= X"01000000";
    when 16#1BBE# => romdata <= X"A20462E0";
    when 16#1BBF# => romdata <= X"C2046004";
    when 16#1BC0# => romdata <= X"82807FFF";
    when 16#1BC1# => romdata <= X"1C800006";
    when 16#1BC2# => romdata <= X"E0046008";
    when 16#1BC3# => romdata <= X"10800026";
    when 16#1BC4# => romdata <= X"D0044000";
    when 16#1BC5# => romdata <= X"0C800023";
    when 16#1BC6# => romdata <= X"A00420CC";
    when 16#1BC7# => romdata <= X"C454200C";
    when 16#1BC8# => romdata <= X"80A0A000";
    when 16#1BC9# => romdata <= X"12BFFFFC";
    when 16#1BCA# => romdata <= X"82807FFF";
    when 16#1BCB# => romdata <= X"82103FFF";
    when 16#1BCC# => romdata <= X"C234200E";
    when 16#1BCD# => romdata <= X"82102001";
    when 16#1BCE# => romdata <= X"C234200C";
    when 16#1BCF# => romdata <= X"A207BFF4";
    when 16#1BD0# => romdata <= X"40000EF5";
    when 16#1BD1# => romdata <= X"90100011";
    when 16#1BD2# => romdata <= X"92102001";
    when 16#1BD3# => romdata <= X"40000F08";
    when 16#1BD4# => romdata <= X"90100011";
    when 16#1BD5# => romdata <= X"92100011";
    when 16#1BD6# => romdata <= X"40000EB6";
    when 16#1BD7# => romdata <= X"90042058";
    when 16#1BD8# => romdata <= X"40000EF8";
    when 16#1BD9# => romdata <= X"90100011";
    when 16#1BDA# => romdata <= X"7FFFFF63";
    when 16#1BDB# => romdata <= X"01000000";
    when 16#1BDC# => romdata <= X"C0240000";
    when 16#1BDD# => romdata <= X"C0242008";
    when 16#1BDE# => romdata <= X"C0242004";
    when 16#1BDF# => romdata <= X"C0242010";
    when 16#1BE0# => romdata <= X"C0242014";
    when 16#1BE1# => romdata <= X"C0242018";
    when 16#1BE2# => romdata <= X"C0242030";
    when 16#1BE3# => romdata <= X"C0242034";
    when 16#1BE4# => romdata <= X"C0242044";
    when 16#1BE5# => romdata <= X"C0242048";
    when 16#1BE6# => romdata <= X"81C7E008";
    when 16#1BE7# => romdata <= X"91E80010";
    when 16#1BE8# => romdata <= X"D0044000";
    when 16#1BE9# => romdata <= X"80A22000";
    when 16#1BEA# => romdata <= X"22800008";
    when 16#1BEB# => romdata <= X"90100018";
    when 16#1BEC# => romdata <= X"10BFFFD3";
    when 16#1BED# => romdata <= X"A2100008";
    when 16#1BEE# => romdata <= X"7FFFFF98";
    when 16#1BEF# => romdata <= X"90100011";
    when 16#1BF0# => romdata <= X"10BFFFCF";
    when 16#1BF1# => romdata <= X"A20462E0";
    when 16#1BF2# => romdata <= X"7FFFFFAF";
    when 16#1BF3# => romdata <= X"92102004";
    when 16#1BF4# => romdata <= X"80A22000";
    when 16#1BF5# => romdata <= X"12BFFFF7";
    when 16#1BF6# => romdata <= X"D0244000";
    when 16#1BF7# => romdata <= X"7FFFFF46";
    when 16#1BF8# => romdata <= X"A0102000";
    when 16#1BF9# => romdata <= X"8210200C";
    when 16#1BFA# => romdata <= X"10BFFFEC";
    when 16#1BFB# => romdata <= X"C2260000";
    when 16#1BFC# => romdata <= X"9DE3BFA0";
    when 16#1BFD# => romdata <= X"7FFFEFE8";
    when 16#1BFE# => romdata <= X"90100018";
    when 16#1BFF# => romdata <= X"21100034";
    when 16#1C00# => romdata <= X"A0142020";
    when 16#1C01# => romdata <= X"C2042008";
    when 16#1C02# => romdata <= X"E2006004";
    when 16#1C03# => romdata <= X"A20C7FFC";
    when 16#1C04# => romdata <= X"82046FEF";
    when 16#1C05# => romdata <= X"B2204019";
    when 16#1C06# => romdata <= X"B20E7000";
    when 16#1C07# => romdata <= X"B2067000";
    when 16#1C08# => romdata <= X"80A66FFF";
    when 16#1C09# => romdata <= X"04800009";
    when 16#1C0A# => romdata <= X"90100018";
    when 16#1C0B# => romdata <= X"7FFFEFE0";
    when 16#1C0C# => romdata <= X"92102000";
    when 16#1C0D# => romdata <= X"C2042008";
    when 16#1C0E# => romdata <= X"82004011";
    when 16#1C0F# => romdata <= X"80A20001";
    when 16#1C10# => romdata <= X"02800007";
    when 16#1C11# => romdata <= X"90100018";
    when 16#1C12# => romdata <= X"90100018";
    when 16#1C13# => romdata <= X"7FFFEFCC";
    when 16#1C14# => romdata <= X"B0102000";
    when 16#1C15# => romdata <= X"81C7E008";
    when 16#1C16# => romdata <= X"81E80000";
    when 16#1C17# => romdata <= X"7FFFEFD4";
    when 16#1C18# => romdata <= X"92200019";
    when 16#1C19# => romdata <= X"80A23FFF";
    when 16#1C1A# => romdata <= X"0280000E";
    when 16#1C1B# => romdata <= X"A2244019";
    when 16#1C1C# => romdata <= X"C4042008";
    when 16#1C1D# => romdata <= X"A2146001";
    when 16#1C1E# => romdata <= X"03100037";
    when 16#1C1F# => romdata <= X"E220A004";
    when 16#1C20# => romdata <= X"90100018";
    when 16#1C21# => romdata <= X"B0102001";
    when 16#1C22# => romdata <= X"C40062FC";
    when 16#1C23# => romdata <= X"B2208019";
    when 16#1C24# => romdata <= X"7FFFEFBB";
    when 16#1C25# => romdata <= X"F22062FC";
    when 16#1C26# => romdata <= X"81C7E008";
    when 16#1C27# => romdata <= X"81E80000";
    when 16#1C28# => romdata <= X"90100018";
    when 16#1C29# => romdata <= X"7FFFEFC2";
    when 16#1C2A# => romdata <= X"92102000";
    when 16#1C2B# => romdata <= X"C2042008";
    when 16#1C2C# => romdata <= X"84220001";
    when 16#1C2D# => romdata <= X"80A0A00F";
    when 16#1C2E# => romdata <= X"04BFFFE4";
    when 16#1C2F# => romdata <= X"07100035";
    when 16#1C30# => romdata <= X"C600E02C";
    when 16#1C31# => romdata <= X"90220003";
    when 16#1C32# => romdata <= X"07100037";
    when 16#1C33# => romdata <= X"8410A001";
    when 16#1C34# => romdata <= X"D020E2FC";
    when 16#1C35# => romdata <= X"10BFFFDD";
    when 16#1C36# => romdata <= X"C4206004";
    when 16#1C37# => romdata <= X"9DE3BFA0";
    when 16#1C38# => romdata <= X"80A66000";
    when 16#1C39# => romdata <= X"02800050";
    when 16#1C3A# => romdata <= X"01000000";
    when 16#1C3B# => romdata <= X"7FFFEFAA";
    when 16#1C3C# => romdata <= X"90100018";
    when 16#1C3D# => romdata <= X"84067FF8";
    when 16#1C3E# => romdata <= X"D800A004";
    when 16#1C3F# => romdata <= X"820B3FFE";
    when 16#1C40# => romdata <= X"09100034";
    when 16#1C41# => romdata <= X"86008001";
    when 16#1C42# => romdata <= X"88112020";
    when 16#1C43# => romdata <= X"DA00E004";
    when 16#1C44# => romdata <= X"D6012008";
    when 16#1C45# => romdata <= X"80A2C003";
    when 16#1C46# => romdata <= X"02800063";
    when 16#1C47# => romdata <= X"9A0B7FFC";
    when 16#1C48# => romdata <= X"DA20E004";
    when 16#1C49# => romdata <= X"808B2001";
    when 16#1C4A# => romdata <= X"1280000E";
    when 16#1C4B# => romdata <= X"98102000";
    when 16#1C4C# => romdata <= X"D8067FF8";
    when 16#1C4D# => romdata <= X"8420800C";
    when 16#1C4E# => romdata <= X"8200400C";
    when 16#1C4F# => romdata <= X"D600A008";
    when 16#1C50# => romdata <= X"98012008";
    when 16#1C51# => romdata <= X"80A2C00C";
    when 16#1C52# => romdata <= X"02800006";
    when 16#1C53# => romdata <= X"98102001";
    when 16#1C54# => romdata <= X"D400A00C";
    when 16#1C55# => romdata <= X"D422E00C";
    when 16#1C56# => romdata <= X"98102000";
    when 16#1C57# => romdata <= X"D622A008";
    when 16#1C58# => romdata <= X"9600C00D";
    when 16#1C59# => romdata <= X"D602E004";
    when 16#1C5A# => romdata <= X"808AE001";
    when 16#1C5B# => romdata <= X"3280000A";
    when 16#1C5C# => romdata <= X"86106001";
    when 16#1C5D# => romdata <= X"80A32000";
    when 16#1C5E# => romdata <= X"0280002D";
    when 16#1C5F# => romdata <= X"8200400D";
    when 16#1C60# => romdata <= X"DA00E008";
    when 16#1C61# => romdata <= X"C600E00C";
    when 16#1C62# => romdata <= X"C623600C";
    when 16#1C63# => romdata <= X"DA20E008";
    when 16#1C64# => romdata <= X"86106001";
    when 16#1C65# => romdata <= X"C2208001";
    when 16#1C66# => romdata <= X"80A32000";
    when 16#1C67# => romdata <= X"12800020";
    when 16#1C68# => romdata <= X"C620A004";
    when 16#1C69# => romdata <= X"80A061FF";
    when 16#1C6A# => romdata <= X"28800030";
    when 16#1C6B# => romdata <= X"83306003";
    when 16#1C6C# => romdata <= X"87306009";
    when 16#1C6D# => romdata <= X"80A0E004";
    when 16#1C6E# => romdata <= X"18800052";
    when 16#1C6F# => romdata <= X"9800E05B";
    when 16#1C70# => romdata <= X"99306006";
    when 16#1C71# => romdata <= X"98032038";
    when 16#1C72# => romdata <= X"9B2B2003";
    when 16#1C73# => romdata <= X"9A01000D";
    when 16#1C74# => romdata <= X"C6036008";
    when 16#1C75# => romdata <= X"80A0C00D";
    when 16#1C76# => romdata <= X"32800008";
    when 16#1C77# => romdata <= X"C800E004";
    when 16#1C78# => romdata <= X"10800052";
    when 16#1C79# => romdata <= X"DA012004";
    when 16#1C7A# => romdata <= X"80A34003";
    when 16#1C7B# => romdata <= X"22800008";
    when 16#1C7C# => romdata <= X"C200E00C";
    when 16#1C7D# => romdata <= X"C800E004";
    when 16#1C7E# => romdata <= X"88093FFC";
    when 16#1C7F# => romdata <= X"80A04004";
    when 16#1C80# => romdata <= X"2ABFFFFA";
    when 16#1C81# => romdata <= X"C600E008";
    when 16#1C82# => romdata <= X"C200E00C";
    when 16#1C83# => romdata <= X"C220A00C";
    when 16#1C84# => romdata <= X"C620A008";
    when 16#1C85# => romdata <= X"C420E00C";
    when 16#1C86# => romdata <= X"C4206008";
    when 16#1C87# => romdata <= X"7FFFEF58";
    when 16#1C88# => romdata <= X"81E80000";
    when 16#1C89# => romdata <= X"81C7E008";
    when 16#1C8A# => romdata <= X"81E80000";
    when 16#1C8B# => romdata <= X"DA00E008";
    when 16#1C8C# => romdata <= X"17100034";
    when 16#1C8D# => romdata <= X"9612E028";
    when 16#1C8E# => romdata <= X"80A3400B";
    when 16#1C8F# => romdata <= X"32BFFFD3";
    when 16#1C90# => romdata <= X"C600E00C";
    when 16#1C91# => romdata <= X"C423600C";
    when 16#1C92# => romdata <= X"C4236008";
    when 16#1C93# => romdata <= X"C2208001";
    when 16#1C94# => romdata <= X"DA20A008";
    when 16#1C95# => romdata <= X"82106001";
    when 16#1C96# => romdata <= X"DA20A00C";
    when 16#1C97# => romdata <= X"C220A004";
    when 16#1C98# => romdata <= X"7FFFEF47";
    when 16#1C99# => romdata <= X"81E80000";
    when 16#1C9A# => romdata <= X"87286003";
    when 16#1C9B# => romdata <= X"86010003";
    when 16#1C9C# => romdata <= X"DA00E008";
    when 16#1C9D# => romdata <= X"C620A00C";
    when 16#1C9E# => romdata <= X"DA20A008";
    when 16#1C9F# => romdata <= X"D8012004";
    when 16#1CA0# => romdata <= X"C423600C";
    when 16#1CA1# => romdata <= X"C420E008";
    when 16#1CA2# => romdata <= X"83386002";
    when 16#1CA3# => romdata <= X"84102001";
    when 16#1CA4# => romdata <= X"83288001";
    when 16#1CA5# => romdata <= X"82130001";
    when 16#1CA6# => romdata <= X"C2212004";
    when 16#1CA7# => romdata <= X"7FFFEF38";
    when 16#1CA8# => romdata <= X"81E80000";
    when 16#1CA9# => romdata <= X"808B2001";
    when 16#1CAA# => romdata <= X"12800009";
    when 16#1CAB# => romdata <= X"82034001";
    when 16#1CAC# => romdata <= X"D8067FF8";
    when 16#1CAD# => romdata <= X"8420800C";
    when 16#1CAE# => romdata <= X"DA00A00C";
    when 16#1CAF# => romdata <= X"C600A008";
    when 16#1CB0# => romdata <= X"8200400C";
    when 16#1CB1# => romdata <= X"C6236008";
    when 16#1CB2# => romdata <= X"DA20E00C";
    when 16#1CB3# => romdata <= X"C4212008";
    when 16#1CB4# => romdata <= X"86106001";
    when 16#1CB5# => romdata <= X"C620A004";
    when 16#1CB6# => romdata <= X"05100035";
    when 16#1CB7# => romdata <= X"C400A028";
    when 16#1CB8# => romdata <= X"80A04002";
    when 16#1CB9# => romdata <= X"0ABFFFCE";
    when 16#1CBA# => romdata <= X"03100037";
    when 16#1CBB# => romdata <= X"D20062F0";
    when 16#1CBC# => romdata <= X"7FFFFF40";
    when 16#1CBD# => romdata <= X"90100018";
    when 16#1CBE# => romdata <= X"7FFFEF21";
    when 16#1CBF# => romdata <= X"81E80000";
    when 16#1CC0# => romdata <= X"80A0E014";
    when 16#1CC1# => romdata <= X"08BFFFB2";
    when 16#1CC2# => romdata <= X"9B2B2003";
    when 16#1CC3# => romdata <= X"80A0E054";
    when 16#1CC4# => romdata <= X"1880000D";
    when 16#1CC5# => romdata <= X"80A0E154";
    when 16#1CC6# => romdata <= X"9930600C";
    when 16#1CC7# => romdata <= X"9803206E";
    when 16#1CC8# => romdata <= X"10BFFFAB";
    when 16#1CC9# => romdata <= X"9B2B2003";
    when 16#1CCA# => romdata <= X"993B2002";
    when 16#1CCB# => romdata <= X"82102001";
    when 16#1CCC# => romdata <= X"8328400C";
    when 16#1CCD# => romdata <= X"82134001";
    when 16#1CCE# => romdata <= X"C2212004";
    when 16#1CCF# => romdata <= X"10BFFFB4";
    when 16#1CD0# => romdata <= X"82100003";
    when 16#1CD1# => romdata <= X"18800006";
    when 16#1CD2# => romdata <= X"80A0E554";
    when 16#1CD3# => romdata <= X"9930600F";
    when 16#1CD4# => romdata <= X"98032077";
    when 16#1CD5# => romdata <= X"10BFFF9E";
    when 16#1CD6# => romdata <= X"9B2B2003";
    when 16#1CD7# => romdata <= X"9A1023F0";
    when 16#1CD8# => romdata <= X"18BFFF9B";
    when 16#1CD9# => romdata <= X"9810207E";
    when 16#1CDA# => romdata <= X"99306012";
    when 16#1CDB# => romdata <= X"9803207C";
    when 16#1CDC# => romdata <= X"10BFFF97";
    when 16#1CDD# => romdata <= X"9B2B2003";
    when 16#1CDE# => romdata <= X"9DE3BFA0";
    when 16#1CDF# => romdata <= X"C2066008";
    when 16#1CE0# => romdata <= X"80A06000";
    when 16#1CE1# => romdata <= X"02800029";
    when 16#1CE2# => romdata <= X"A0100018";
    when 16#1CE3# => romdata <= X"C416200C";
    when 16#1CE4# => romdata <= X"8088A008";
    when 16#1CE5# => romdata <= X"028000F3";
    when 16#1CE6# => romdata <= X"82100002";
    when 16#1CE7# => romdata <= X"C6062010";
    when 16#1CE8# => romdata <= X"80A0E000";
    when 16#1CE9# => romdata <= X"028000F0";
    when 16#1CEA# => romdata <= X"90100010";
    when 16#1CEB# => romdata <= X"8088A002";
    when 16#1CEC# => romdata <= X"E2064000";
    when 16#1CED# => romdata <= X"A6102000";
    when 16#1CEE# => romdata <= X"0280001F";
    when 16#1CEF# => romdata <= X"A4102000";
    when 16#1CF0# => romdata <= X"80A4A000";
    when 16#1CF1# => romdata <= X"02800015";
    when 16#1CF2# => romdata <= X"92100013";
    when 16#1CF3# => romdata <= X"80A4A400";
    when 16#1CF4# => romdata <= X"08800003";
    when 16#1CF5# => romdata <= X"94100012";
    when 16#1CF6# => romdata <= X"94102400";
    when 16#1CF7# => romdata <= X"C2042024";
    when 16#1CF8# => romdata <= X"9FC04000";
    when 16#1CF9# => romdata <= X"D004201C";
    when 16#1CFA# => romdata <= X"80A22000";
    when 16#1CFB# => romdata <= X"04800098";
    when 16#1CFC# => romdata <= X"A4248008";
    when 16#1CFD# => romdata <= X"C2066008";
    when 16#1CFE# => romdata <= X"82204008";
    when 16#1CFF# => romdata <= X"80A06000";
    when 16#1D00# => romdata <= X"0280000A";
    when 16#1D01# => romdata <= X"C2266008";
    when 16#1D02# => romdata <= X"A604C008";
    when 16#1D03# => romdata <= X"80A4A000";
    when 16#1D04# => romdata <= X"12BFFFEF";
    when 16#1D05# => romdata <= X"92100013";
    when 16#1D06# => romdata <= X"E6044000";
    when 16#1D07# => romdata <= X"E4046004";
    when 16#1D08# => romdata <= X"10BFFFE8";
    when 16#1D09# => romdata <= X"A2046008";
    when 16#1D0A# => romdata <= X"B0102000";
    when 16#1D0B# => romdata <= X"81C7E008";
    when 16#1D0C# => romdata <= X"81E80000";
    when 16#1D0D# => romdata <= X"2D100032";
    when 16#1D0E# => romdata <= X"8088A001";
    when 16#1D0F# => romdata <= X"AC15A2C8";
    when 16#1D10# => romdata <= X"0280004E";
    when 16#1D11# => romdata <= X"A8102000";
    when 16#1D12# => romdata <= X"AE102000";
    when 16#1D13# => romdata <= X"AC102000";
    when 16#1D14# => romdata <= X"A6102000";
    when 16#1D15# => romdata <= X"80A4E000";
    when 16#1D16# => romdata <= X"2280002B";
    when 16#1D17# => romdata <= X"EC044000";
    when 16#1D18# => romdata <= X"80A5E000";
    when 16#1D19# => romdata <= X"028000B5";
    when 16#1D1A# => romdata <= X"90100016";
    when 16#1D1B# => romdata <= X"80A50013";
    when 16#1D1C# => romdata <= X"08800003";
    when 16#1D1D# => romdata <= X"AA100014";
    when 16#1D1E# => romdata <= X"AA100013";
    when 16#1D1F# => romdata <= X"D4042014";
    when 16#1D20# => romdata <= X"E4042008";
    when 16#1D21# => romdata <= X"A4028012";
    when 16#1D22# => romdata <= X"80A54012";
    when 16#1D23# => romdata <= X"0480008D";
    when 16#1D24# => romdata <= X"D0040000";
    when 16#1D25# => romdata <= X"C2042010";
    when 16#1D26# => romdata <= X"80A20001";
    when 16#1D27# => romdata <= X"0880008A";
    when 16#1D28# => romdata <= X"80A5400A";
    when 16#1D29# => romdata <= X"92100016";
    when 16#1D2A# => romdata <= X"4000022C";
    when 16#1D2B# => romdata <= X"94100012";
    when 16#1D2C# => romdata <= X"C2040000";
    when 16#1D2D# => romdata <= X"82004012";
    when 16#1D2E# => romdata <= X"C2240000";
    when 16#1D2F# => romdata <= X"7FFFFDA2";
    when 16#1D30# => romdata <= X"90100010";
    when 16#1D31# => romdata <= X"80A22000";
    when 16#1D32# => romdata <= X"32800062";
    when 16#1D33# => romdata <= X"C214200C";
    when 16#1D34# => romdata <= X"A8A50012";
    when 16#1D35# => romdata <= X"02800088";
    when 16#1D36# => romdata <= X"01000000";
    when 16#1D37# => romdata <= X"C2066008";
    when 16#1D38# => romdata <= X"82204012";
    when 16#1D39# => romdata <= X"80A06000";
    when 16#1D3A# => romdata <= X"02BFFFD0";
    when 16#1D3B# => romdata <= X"C2266008";
    when 16#1D3C# => romdata <= X"A624C012";
    when 16#1D3D# => romdata <= X"80A4E000";
    when 16#1D3E# => romdata <= X"12BFFFDA";
    when 16#1D3F# => romdata <= X"AC058012";
    when 16#1D40# => romdata <= X"EC044000";
    when 16#1D41# => romdata <= X"E6046004";
    when 16#1D42# => romdata <= X"AE102000";
    when 16#1D43# => romdata <= X"10BFFFD2";
    when 16#1D44# => romdata <= X"A2046008";
    when 16#1D45# => romdata <= X"D0040000";
    when 16#1D46# => romdata <= X"80A48015";
    when 16#1D47# => romdata <= X"1A800005";
    when 16#1D48# => romdata <= X"94100015";
    when 16#1D49# => romdata <= X"AA100012";
    when 16#1D4A# => romdata <= X"A6100012";
    when 16#1D4B# => romdata <= X"94100015";
    when 16#1D4C# => romdata <= X"4000020A";
    when 16#1D4D# => romdata <= X"92100014";
    when 16#1D4E# => romdata <= X"C4042008";
    when 16#1D4F# => romdata <= X"C2040000";
    when 16#1D50# => romdata <= X"A6208013";
    when 16#1D51# => romdata <= X"AA004015";
    when 16#1D52# => romdata <= X"E6242008";
    when 16#1D53# => romdata <= X"EA240000";
    when 16#1D54# => romdata <= X"A6100012";
    when 16#1D55# => romdata <= X"AA100012";
    when 16#1D56# => romdata <= X"C2066008";
    when 16#1D57# => romdata <= X"A6204013";
    when 16#1D58# => romdata <= X"80A4E000";
    when 16#1D59# => romdata <= X"02BFFFB1";
    when 16#1D5A# => romdata <= X"E6266008";
    when 16#1D5B# => romdata <= X"C214200C";
    when 16#1D5C# => romdata <= X"A4248015";
    when 16#1D5D# => romdata <= X"A8050015";
    when 16#1D5E# => romdata <= X"80A4A000";
    when 16#1D5F# => romdata <= X"2280001E";
    when 16#1D60# => romdata <= X"E8044000";
    when 16#1D61# => romdata <= X"83286010";
    when 16#1D62# => romdata <= X"83306010";
    when 16#1D63# => romdata <= X"80886200";
    when 16#1D64# => romdata <= X"0280001C";
    when 16#1D65# => romdata <= X"E6042008";
    when 16#1D66# => romdata <= X"80A48013";
    when 16#1D67# => romdata <= X"08BFFFDE";
    when 16#1D68# => romdata <= X"AA100013";
    when 16#1D69# => romdata <= X"80886080";
    when 16#1D6A# => romdata <= X"22BFFFDC";
    when 16#1D6B# => romdata <= X"D0040000";
    when 16#1D6C# => romdata <= X"D2042010";
    when 16#1D6D# => romdata <= X"EA040000";
    when 16#1D6E# => romdata <= X"D0058000";
    when 16#1D6F# => romdata <= X"AA254009";
    when 16#1D70# => romdata <= X"A6048015";
    when 16#1D71# => romdata <= X"4000060C";
    when 16#1D72# => romdata <= X"94100013";
    when 16#1D73# => romdata <= X"82922000";
    when 16#1D74# => romdata <= X"0280006D";
    when 16#1D75# => romdata <= X"90004015";
    when 16#1D76# => romdata <= X"E6242014";
    when 16#1D77# => romdata <= X"C2242010";
    when 16#1D78# => romdata <= X"D0240000";
    when 16#1D79# => romdata <= X"E4242008";
    when 16#1D7A# => romdata <= X"A6100012";
    when 16#1D7B# => romdata <= X"10BFFFCB";
    when 16#1D7C# => romdata <= X"AA100012";
    when 16#1D7D# => romdata <= X"E4046004";
    when 16#1D7E# => romdata <= X"10BFFFE0";
    when 16#1D7F# => romdata <= X"A2046008";
    when 16#1D80# => romdata <= X"80A4C012";
    when 16#1D81# => romdata <= X"D0040000";
    when 16#1D82# => romdata <= X"1A800016";
    when 16#1D83# => romdata <= X"AA100013";
    when 16#1D84# => romdata <= X"C2042010";
    when 16#1D85# => romdata <= X"80A20001";
    when 16#1D86# => romdata <= X"28800013";
    when 16#1D87# => romdata <= X"D4042014";
    when 16#1D88# => romdata <= X"92100014";
    when 16#1D89# => romdata <= X"400001CD";
    when 16#1D8A# => romdata <= X"94100013";
    when 16#1D8B# => romdata <= X"C2040000";
    when 16#1D8C# => romdata <= X"82004013";
    when 16#1D8D# => romdata <= X"C2240000";
    when 16#1D8E# => romdata <= X"7FFFFD43";
    when 16#1D8F# => romdata <= X"90100010";
    when 16#1D90# => romdata <= X"80A22000";
    when 16#1D91# => romdata <= X"22BFFFC6";
    when 16#1D92# => romdata <= X"C2066008";
    when 16#1D93# => romdata <= X"C214200C";
    when 16#1D94# => romdata <= X"82106040";
    when 16#1D95# => romdata <= X"C234200C";
    when 16#1D96# => romdata <= X"81C7E008";
    when 16#1D97# => romdata <= X"91E83FFF";
    when 16#1D98# => romdata <= X"D4042014";
    when 16#1D99# => romdata <= X"80A4800A";
    when 16#1D9A# => romdata <= X"0A80000B";
    when 16#1D9B# => romdata <= X"92100014";
    when 16#1D9C# => romdata <= X"C2042024";
    when 16#1D9D# => romdata <= X"D004201C";
    when 16#1D9E# => romdata <= X"9FC04000";
    when 16#1D9F# => romdata <= X"92100014";
    when 16#1DA0# => romdata <= X"A6922000";
    when 16#1DA1# => romdata <= X"24BFFFF3";
    when 16#1DA2# => romdata <= X"C214200C";
    when 16#1DA3# => romdata <= X"10BFFFB3";
    when 16#1DA4# => romdata <= X"AA100013";
    when 16#1DA5# => romdata <= X"400001B1";
    when 16#1DA6# => romdata <= X"94100012";
    when 16#1DA7# => romdata <= X"C4042008";
    when 16#1DA8# => romdata <= X"C2040000";
    when 16#1DA9# => romdata <= X"84208012";
    when 16#1DAA# => romdata <= X"82004012";
    when 16#1DAB# => romdata <= X"C4242008";
    when 16#1DAC# => romdata <= X"C2240000";
    when 16#1DAD# => romdata <= X"A6100012";
    when 16#1DAE# => romdata <= X"10BFFFA8";
    when 16#1DAF# => romdata <= X"AA100012";
    when 16#1DB0# => romdata <= X"80A5400A";
    when 16#1DB1# => romdata <= X"06800013";
    when 16#1DB2# => romdata <= X"92100016";
    when 16#1DB3# => romdata <= X"C2042024";
    when 16#1DB4# => romdata <= X"D004201C";
    when 16#1DB5# => romdata <= X"9FC04000";
    when 16#1DB6# => romdata <= X"92100016";
    when 16#1DB7# => romdata <= X"A4922000";
    when 16#1DB8# => romdata <= X"24BFFFDC";
    when 16#1DB9# => romdata <= X"C214200C";
    when 16#1DBA# => romdata <= X"A8A50012";
    when 16#1DBB# => romdata <= X"32BFFF7D";
    when 16#1DBC# => romdata <= X"C2066008";
    when 16#1DBD# => romdata <= X"7FFFFD14";
    when 16#1DBE# => romdata <= X"90100010";
    when 16#1DBF# => romdata <= X"80A22000";
    when 16#1DC0# => romdata <= X"12BFFFD3";
    when 16#1DC1# => romdata <= X"AE102000";
    when 16#1DC2# => romdata <= X"10BFFF76";
    when 16#1DC3# => romdata <= X"C2066008";
    when 16#1DC4# => romdata <= X"40000192";
    when 16#1DC5# => romdata <= X"94100015";
    when 16#1DC6# => romdata <= X"C4042008";
    when 16#1DC7# => romdata <= X"C2040000";
    when 16#1DC8# => romdata <= X"84208015";
    when 16#1DC9# => romdata <= X"82004015";
    when 16#1DCA# => romdata <= X"C4242008";
    when 16#1DCB# => romdata <= X"C2240000";
    when 16#1DCC# => romdata <= X"10BFFF68";
    when 16#1DCD# => romdata <= X"A4100015";
    when 16#1DCE# => romdata <= X"9210200A";
    when 16#1DCF# => romdata <= X"94100013";
    when 16#1DD0# => romdata <= X"4000010B";
    when 16#1DD1# => romdata <= X"A804E001";
    when 16#1DD2# => romdata <= X"80A22000";
    when 16#1DD3# => romdata <= X"02BFFF48";
    when 16#1DD4# => romdata <= X"AE102001";
    when 16#1DD5# => romdata <= X"A8022001";
    when 16#1DD6# => romdata <= X"10BFFF45";
    when 16#1DD7# => romdata <= X"A8250016";
    when 16#1DD8# => romdata <= X"90100010";
    when 16#1DD9# => romdata <= X"7FFFF764";
    when 16#1DDA# => romdata <= X"B0103FFF";
    when 16#1DDB# => romdata <= X"80A22000";
    when 16#1DDC# => romdata <= X"12BFFF2F";
    when 16#1DDD# => romdata <= X"01000000";
    when 16#1DDE# => romdata <= X"C214200C";
    when 16#1DDF# => romdata <= X"10BFFF0C";
    when 16#1DE0# => romdata <= X"84100001";
    when 16#1DE1# => romdata <= X"D0058000";
    when 16#1DE2# => romdata <= X"7FFFFE55";
    when 16#1DE3# => romdata <= X"D2042010";
    when 16#1DE4# => romdata <= X"10BFFFB0";
    when 16#1DE5# => romdata <= X"C214200C";
    when 16#1DE6# => romdata <= X"9DE3BFA0";
    when 16#1DE7# => romdata <= X"7FFFFD6E";
    when 16#1DE8# => romdata <= X"A0100018";
    when 16#1DE9# => romdata <= X"A68422E0";
    when 16#1DEA# => romdata <= X"02800031";
    when 16#1DEB# => romdata <= X"B0102000";
    when 16#1DEC# => romdata <= X"E404E004";
    when 16#1DED# => romdata <= X"A484BFFF";
    when 16#1DEE# => romdata <= X"1C800014";
    when 16#1DEF# => romdata <= X"E204E008";
    when 16#1DF0# => romdata <= X"10800028";
    when 16#1DF1# => romdata <= X"E604C000";
    when 16#1DF2# => romdata <= X"C454600E";
    when 16#1DF3# => romdata <= X"92100011";
    when 16#1DF4# => romdata <= X"80A0BFFF";
    when 16#1DF5# => romdata <= X"02800006";
    when 16#1DF6# => romdata <= X"90100010";
    when 16#1DF7# => romdata <= X"9FC64000";
    when 16#1DF8# => romdata <= X"01000000";
    when 16#1DF9# => romdata <= X"C214600C";
    when 16#1DFA# => romdata <= X"B0160008";
    when 16#1DFB# => romdata <= X"80886200";
    when 16#1DFC# => romdata <= X"02800016";
    when 16#1DFD# => romdata <= X"A8046058";
    when 16#1DFE# => romdata <= X"A484BFFF";
    when 16#1DFF# => romdata <= X"2C800019";
    when 16#1E00# => romdata <= X"E604C000";
    when 16#1E01# => romdata <= X"A20460CC";
    when 16#1E02# => romdata <= X"C214600C";
    when 16#1E03# => romdata <= X"85286010";
    when 16#1E04# => romdata <= X"80A0A000";
    when 16#1E05# => romdata <= X"22BFFFFA";
    when 16#1E06# => romdata <= X"A484BFFF";
    when 16#1E07# => romdata <= X"8530A010";
    when 16#1E08# => romdata <= X"8088A200";
    when 16#1E09# => romdata <= X"32BFFFEA";
    when 16#1E0A# => romdata <= X"C454600E";
    when 16#1E0B# => romdata <= X"A8046058";
    when 16#1E0C# => romdata <= X"40000C98";
    when 16#1E0D# => romdata <= X"90100014";
    when 16#1E0E# => romdata <= X"C254600C";
    when 16#1E0F# => romdata <= X"80A06000";
    when 16#1E10# => romdata <= X"12BFFFE2";
    when 16#1E11# => romdata <= X"C214600C";
    when 16#1E12# => romdata <= X"40000CA8";
    when 16#1E13# => romdata <= X"90100014";
    when 16#1E14# => romdata <= X"A484BFFF";
    when 16#1E15# => romdata <= X"3CBFFFED";
    when 16#1E16# => romdata <= X"A20460CC";
    when 16#1E17# => romdata <= X"E604C000";
    when 16#1E18# => romdata <= X"80A4E000";
    when 16#1E19# => romdata <= X"32BFFFD4";
    when 16#1E1A# => romdata <= X"E404E004";
    when 16#1E1B# => romdata <= X"7FFFFD22";
    when 16#1E1C# => romdata <= X"01000000";
    when 16#1E1D# => romdata <= X"81C7E008";
    when 16#1E1E# => romdata <= X"81E80000";
    when 16#1E1F# => romdata <= X"9DE3BFA0";
    when 16#1E20# => romdata <= X"7FFFFD35";
    when 16#1E21# => romdata <= X"01000000";
    when 16#1E22# => romdata <= X"A48622E0";
    when 16#1E23# => romdata <= X"02800030";
    when 16#1E24# => romdata <= X"B0102000";
    when 16#1E25# => romdata <= X"E204A004";
    when 16#1E26# => romdata <= X"A2847FFF";
    when 16#1E27# => romdata <= X"1C800013";
    when 16#1E28# => romdata <= X"E004A008";
    when 16#1E29# => romdata <= X"10800027";
    when 16#1E2A# => romdata <= X"E4048000";
    when 16#1E2B# => romdata <= X"C454200E";
    when 16#1E2C# => romdata <= X"80A0BFFF";
    when 16#1E2D# => romdata <= X"02800006";
    when 16#1E2E# => romdata <= X"90100010";
    when 16#1E2F# => romdata <= X"9FC64000";
    when 16#1E30# => romdata <= X"01000000";
    when 16#1E31# => romdata <= X"C214200C";
    when 16#1E32# => romdata <= X"B0160008";
    when 16#1E33# => romdata <= X"80886200";
    when 16#1E34# => romdata <= X"02800016";
    when 16#1E35# => romdata <= X"A6042058";
    when 16#1E36# => romdata <= X"A2847FFF";
    when 16#1E37# => romdata <= X"2C800019";
    when 16#1E38# => romdata <= X"E4048000";
    when 16#1E39# => romdata <= X"A00420CC";
    when 16#1E3A# => romdata <= X"C214200C";
    when 16#1E3B# => romdata <= X"85286010";
    when 16#1E3C# => romdata <= X"80A0A000";
    when 16#1E3D# => romdata <= X"22BFFFFA";
    when 16#1E3E# => romdata <= X"A2847FFF";
    when 16#1E3F# => romdata <= X"8530A010";
    when 16#1E40# => romdata <= X"8088A200";
    when 16#1E41# => romdata <= X"32BFFFEB";
    when 16#1E42# => romdata <= X"C454200E";
    when 16#1E43# => romdata <= X"A6042058";
    when 16#1E44# => romdata <= X"40000C60";
    when 16#1E45# => romdata <= X"90100013";
    when 16#1E46# => romdata <= X"C254200C";
    when 16#1E47# => romdata <= X"80A06000";
    when 16#1E48# => romdata <= X"12BFFFE3";
    when 16#1E49# => romdata <= X"C214200C";
    when 16#1E4A# => romdata <= X"40000C70";
    when 16#1E4B# => romdata <= X"90100013";
    when 16#1E4C# => romdata <= X"A2847FFF";
    when 16#1E4D# => romdata <= X"3CBFFFED";
    when 16#1E4E# => romdata <= X"A00420CC";
    when 16#1E4F# => romdata <= X"E4048000";
    when 16#1E50# => romdata <= X"80A4A000";
    when 16#1E51# => romdata <= X"32BFFFD5";
    when 16#1E52# => romdata <= X"E204A004";
    when 16#1E53# => romdata <= X"7FFFFCEA";
    when 16#1E54# => romdata <= X"01000000";
    when 16#1E55# => romdata <= X"81C7E008";
    when 16#1E56# => romdata <= X"81E80000";
    when 16#1E57# => romdata <= X"03100032";
    when 16#1E58# => romdata <= X"81C3E008";
    when 16#1E59# => romdata <= X"D0006148";
    when 16#1E5A# => romdata <= X"11100032";
    when 16#1E5B# => romdata <= X"81C3E008";
    when 16#1E5C# => romdata <= X"90122118";
    when 16#1E5D# => romdata <= X"11100032";
    when 16#1E5E# => romdata <= X"81C3E008";
    when 16#1E5F# => romdata <= X"90122118";
    when 16#1E60# => romdata <= X"9DE3BFA0";
    when 16#1E61# => romdata <= X"A0100018";
    when 16#1E62# => romdata <= X"80A6A000";
    when 16#1E63# => romdata <= X"31100032";
    when 16#1E64# => romdata <= X"02800014";
    when 16#1E65# => romdata <= X"B0162000";
    when 16#1E66# => romdata <= X"9010001A";
    when 16#1E67# => romdata <= X"92100018";
    when 16#1E68# => romdata <= X"7FFFEB05";
    when 16#1E69# => romdata <= X"23100032";
    when 16#1E6A# => romdata <= X"80A22000";
    when 16#1E6B# => romdata <= X"12800006";
    when 16#1E6C# => romdata <= X"9010001A";
    when 16#1E6D# => romdata <= X"F4242034";
    when 16#1E6E# => romdata <= X"F2242030";
    when 16#1E6F# => romdata <= X"81C7E008";
    when 16#1E70# => romdata <= X"91EC6000";
    when 16#1E71# => romdata <= X"13100031";
    when 16#1E72# => romdata <= X"B0102000";
    when 16#1E73# => romdata <= X"7FFFEAFA";
    when 16#1E74# => romdata <= X"92126100";
    when 16#1E75# => romdata <= X"80A22000";
    when 16#1E76# => romdata <= X"22BFFFF8";
    when 16#1E77# => romdata <= X"F4242034";
    when 16#1E78# => romdata <= X"81C7E008";
    when 16#1E79# => romdata <= X"81E80000";
    when 16#1E7A# => romdata <= X"82100008";
    when 16#1E7B# => romdata <= X"05100032";
    when 16#1E7C# => romdata <= X"D000A2C8";
    when 16#1E7D# => romdata <= X"94100009";
    when 16#1E7E# => romdata <= X"92100001";
    when 16#1E7F# => romdata <= X"8213C000";
    when 16#1E80# => romdata <= X"7FFFFFE0";
    when 16#1E81# => romdata <= X"9E104000";
    when 16#1E82# => romdata <= X"01000000";
    when 16#1E83# => romdata <= X"9DE3BF60";
    when 16#1E84# => romdata <= X"C216200C";
    when 16#1E85# => romdata <= X"80886002";
    when 16#1E86# => romdata <= X"3280003B";
    when 16#1E87# => romdata <= X"82062043";
    when 16#1E88# => romdata <= X"D256200E";
    when 16#1E89# => romdata <= X"80A26000";
    when 16#1E8A# => romdata <= X"06800017";
    when 16#1E8B# => romdata <= X"21100032";
    when 16#1E8C# => romdata <= X"D00422C8";
    when 16#1E8D# => romdata <= X"400007CC";
    when 16#1E8E# => romdata <= X"9407BFC0";
    when 16#1E8F# => romdata <= X"80A22000";
    when 16#1E90# => romdata <= X"06800010";
    when 16#1E91# => romdata <= X"C417BFC8";
    when 16#1E92# => romdata <= X"0300003C";
    when 16#1E93# => romdata <= X"82088001";
    when 16#1E94# => romdata <= X"05000008";
    when 16#1E95# => romdata <= X"84184002";
    when 16#1E96# => romdata <= X"80A00002";
    when 16#1E97# => romdata <= X"05000020";
    when 16#1E98# => romdata <= X"A2603FFF";
    when 16#1E99# => romdata <= X"80A04002";
    when 16#1E9A# => romdata <= X"2280002D";
    when 16#1E9B# => romdata <= X"C4062028";
    when 16#1E9C# => romdata <= X"C216200C";
    when 16#1E9D# => romdata <= X"82106800";
    when 16#1E9E# => romdata <= X"10800006";
    when 16#1E9F# => romdata <= X"C236200C";
    when 16#1EA0# => romdata <= X"C216200C";
    when 16#1EA1# => romdata <= X"82106800";
    when 16#1EA2# => romdata <= X"A2102000";
    when 16#1EA3# => romdata <= X"C236200C";
    when 16#1EA4# => romdata <= X"D00422C8";
    when 16#1EA5# => romdata <= X"7FFFEB84";
    when 16#1EA6# => romdata <= X"92102400";
    when 16#1EA7# => romdata <= X"80A22000";
    when 16#1EA8# => romdata <= X"02800029";
    when 16#1EA9# => romdata <= X"03100032";
    when 16#1EAA# => romdata <= X"C416200C";
    when 16#1EAB# => romdata <= X"C20062C8";
    when 16#1EAC# => romdata <= X"8410A080";
    when 16#1EAD# => romdata <= X"D0262010";
    when 16#1EAE# => romdata <= X"D0260000";
    when 16#1EAF# => romdata <= X"C436200C";
    when 16#1EB0# => romdata <= X"0510001B";
    when 16#1EB1# => romdata <= X"8410A0A0";
    when 16#1EB2# => romdata <= X"C420603C";
    when 16#1EB3# => romdata <= X"82102400";
    when 16#1EB4# => romdata <= X"80A46000";
    when 16#1EB5# => romdata <= X"0280000A";
    when 16#1EB6# => romdata <= X"C2262014";
    when 16#1EB7# => romdata <= X"40000970";
    when 16#1EB8# => romdata <= X"D056200E";
    when 16#1EB9# => romdata <= X"80A22000";
    when 16#1EBA# => romdata <= X"0280001F";
    when 16#1EBB# => romdata <= X"01000000";
    when 16#1EBC# => romdata <= X"C216200C";
    when 16#1EBD# => romdata <= X"82106001";
    when 16#1EBE# => romdata <= X"C236200C";
    when 16#1EBF# => romdata <= X"81C7E008";
    when 16#1EC0# => romdata <= X"81E80000";
    when 16#1EC1# => romdata <= X"C2262010";
    when 16#1EC2# => romdata <= X"C2260000";
    when 16#1EC3# => romdata <= X"82102001";
    when 16#1EC4# => romdata <= X"C2262014";
    when 16#1EC5# => romdata <= X"81C7E008";
    when 16#1EC6# => romdata <= X"81E80000";
    when 16#1EC7# => romdata <= X"03100025";
    when 16#1EC8# => romdata <= X"8210611C";
    when 16#1EC9# => romdata <= X"80A08001";
    when 16#1ECA# => romdata <= X"12BFFFD3";
    when 16#1ECB# => romdata <= X"C216200C";
    when 16#1ECC# => romdata <= X"82106400";
    when 16#1ECD# => romdata <= X"84102400";
    when 16#1ECE# => romdata <= X"C426204C";
    when 16#1ECF# => romdata <= X"10BFFFD5";
    when 16#1ED0# => romdata <= X"C236200C";
    when 16#1ED1# => romdata <= X"C416200C";
    when 16#1ED2# => romdata <= X"8410A002";
    when 16#1ED3# => romdata <= X"82062043";
    when 16#1ED4# => romdata <= X"C2262010";
    when 16#1ED5# => romdata <= X"C2260000";
    when 16#1ED6# => romdata <= X"C436200C";
    when 16#1ED7# => romdata <= X"82102001";
    when 16#1ED8# => romdata <= X"C2262014";
    when 16#1ED9# => romdata <= X"81C7E008";
    when 16#1EDA# => romdata <= X"81E80000";
    when 16#1EDB# => romdata <= X"9DE3BFA0";
    when 16#1EDC# => romdata <= X"B20E60FF";
    when 16#1EDD# => romdata <= X"80A6A003";
    when 16#1EDE# => romdata <= X"08800029";
    when 16#1EDF# => romdata <= X"82100018";
    when 16#1EE0# => romdata <= X"808E2003";
    when 16#1EE1# => romdata <= X"1280002E";
    when 16#1EE2# => romdata <= X"9B2E6008";
    when 16#1EE3# => romdata <= X"093FBFBF";
    when 16#1EE4# => romdata <= X"9A034019";
    when 16#1EE5# => romdata <= X"07202020";
    when 16#1EE6# => romdata <= X"9B2B6008";
    when 16#1EE7# => romdata <= X"881122FF";
    when 16#1EE8# => romdata <= X"9A034019";
    when 16#1EE9# => romdata <= X"8610E080";
    when 16#1EEA# => romdata <= X"9B2B6008";
    when 16#1EEB# => romdata <= X"9A034019";
    when 16#1EEC# => romdata <= X"C2060000";
    when 16#1EED# => romdata <= X"821B4001";
    when 16#1EEE# => romdata <= X"84004004";
    when 16#1EEF# => romdata <= X"82288001";
    when 16#1EF0# => romdata <= X"80884003";
    when 16#1EF1# => romdata <= X"02800012";
    when 16#1EF2# => romdata <= X"B406BFFC";
    when 16#1EF3# => romdata <= X"C20E0000";
    when 16#1EF4# => romdata <= X"80A04019";
    when 16#1EF5# => romdata <= X"02800020";
    when 16#1EF6# => romdata <= X"01000000";
    when 16#1EF7# => romdata <= X"C20E2001";
    when 16#1EF8# => romdata <= X"80A04019";
    when 16#1EF9# => romdata <= X"0280001A";
    when 16#1EFA# => romdata <= X"82062001";
    when 16#1EFB# => romdata <= X"C20E2002";
    when 16#1EFC# => romdata <= X"80A04019";
    when 16#1EFD# => romdata <= X"02800016";
    when 16#1EFE# => romdata <= X"82062002";
    when 16#1EFF# => romdata <= X"C20E2003";
    when 16#1F00# => romdata <= X"80A04019";
    when 16#1F01# => romdata <= X"02800012";
    when 16#1F02# => romdata <= X"82062003";
    when 16#1F03# => romdata <= X"80A6A003";
    when 16#1F04# => romdata <= X"18BFFFE8";
    when 16#1F05# => romdata <= X"B0062004";
    when 16#1F06# => romdata <= X"82100018";
    when 16#1F07# => romdata <= X"80A6A000";
    when 16#1F08# => romdata <= X"32800008";
    when 16#1F09# => romdata <= X"C4084000";
    when 16#1F0A# => romdata <= X"81C7E008";
    when 16#1F0B# => romdata <= X"91E82000";
    when 16#1F0C# => romdata <= X"80A6A000";
    when 16#1F0D# => romdata <= X"02BFFFFD";
    when 16#1F0E# => romdata <= X"82006001";
    when 16#1F0F# => romdata <= X"C4084000";
    when 16#1F10# => romdata <= X"80A08019";
    when 16#1F11# => romdata <= X"12BFFFFB";
    when 16#1F12# => romdata <= X"B406BFFF";
    when 16#1F13# => romdata <= X"81C7E008";
    when 16#1F14# => romdata <= X"91E80001";
    when 16#1F15# => romdata <= X"81C7E008";
    when 16#1F16# => romdata <= X"81E80000";
    when 16#1F17# => romdata <= X"9DE3BFA0";
    when 16#1F18# => romdata <= X"80A6A00F";
    when 16#1F19# => romdata <= X"9A100018";
    when 16#1F1A# => romdata <= X"88100019";
    when 16#1F1B# => romdata <= X"08800006";
    when 16#1F1C# => romdata <= X"8610001A";
    when 16#1F1D# => romdata <= X"82164018";
    when 16#1F1E# => romdata <= X"80886003";
    when 16#1F1F# => romdata <= X"0280000D";
    when 16#1F20# => romdata <= X"84100019";
    when 16#1F21# => romdata <= X"80A0E000";
    when 16#1F22# => romdata <= X"02800008";
    when 16#1F23# => romdata <= X"82102000";
    when 16#1F24# => romdata <= X"C4090001";
    when 16#1F25# => romdata <= X"C42B4001";
    when 16#1F26# => romdata <= X"82006001";
    when 16#1F27# => romdata <= X"80A04003";
    when 16#1F28# => romdata <= X"32BFFFFD";
    when 16#1F29# => romdata <= X"C4090001";
    when 16#1F2A# => romdata <= X"81C7E008";
    when 16#1F2B# => romdata <= X"81E80000";
    when 16#1F2C# => romdata <= X"82100018";
    when 16#1F2D# => romdata <= X"DA008000";
    when 16#1F2E# => romdata <= X"DA204000";
    when 16#1F2F# => romdata <= X"8600FFF0";
    when 16#1F30# => romdata <= X"80A0E00F";
    when 16#1F31# => romdata <= X"DA00A004";
    when 16#1F32# => romdata <= X"DA206004";
    when 16#1F33# => romdata <= X"DA00A008";
    when 16#1F34# => romdata <= X"DA206008";
    when 16#1F35# => romdata <= X"DA00A00C";
    when 16#1F36# => romdata <= X"DA20600C";
    when 16#1F37# => romdata <= X"8400A010";
    when 16#1F38# => romdata <= X"18BFFFF5";
    when 16#1F39# => romdata <= X"82006010";
    when 16#1F3A# => romdata <= X"B406BFF0";
    when 16#1F3B# => romdata <= X"9B36A004";
    when 16#1F3C# => romdata <= X"832B6004";
    when 16#1F3D# => romdata <= X"9A036001";
    when 16#1F3E# => romdata <= X"B4268001";
    when 16#1F3F# => romdata <= X"9B2B6004";
    when 16#1F40# => romdata <= X"80A6A003";
    when 16#1F41# => romdata <= X"8806400D";
    when 16#1F42# => romdata <= X"8610001A";
    when 16#1F43# => romdata <= X"08BFFFDE";
    when 16#1F44# => romdata <= X"9A06000D";
    when 16#1F45# => romdata <= X"82102000";
    when 16#1F46# => romdata <= X"C4010001";
    when 16#1F47# => romdata <= X"C4234001";
    when 16#1F48# => romdata <= X"82006004";
    when 16#1F49# => romdata <= X"84268001";
    when 16#1F4A# => romdata <= X"80A0A003";
    when 16#1F4B# => romdata <= X"38BFFFFC";
    when 16#1F4C# => romdata <= X"C4010001";
    when 16#1F4D# => romdata <= X"B406BFFC";
    when 16#1F4E# => romdata <= X"8336A002";
    when 16#1F4F# => romdata <= X"87286002";
    when 16#1F50# => romdata <= X"82006001";
    when 16#1F51# => romdata <= X"86268003";
    when 16#1F52# => romdata <= X"83286002";
    when 16#1F53# => romdata <= X"88010001";
    when 16#1F54# => romdata <= X"10BFFFCD";
    when 16#1F55# => romdata <= X"9A034001";
    when 16#1F56# => romdata <= X"9DE3BFA0";
    when 16#1F57# => romdata <= X"80A60019";
    when 16#1F58# => romdata <= X"9A100018";
    when 16#1F59# => romdata <= X"88100019";
    when 16#1F5A# => romdata <= X"08800013";
    when 16#1F5B# => romdata <= X"8610001A";
    when 16#1F5C# => romdata <= X"8206401A";
    when 16#1F5D# => romdata <= X"80A60001";
    when 16#1F5E# => romdata <= X"1A800010";
    when 16#1F5F# => romdata <= X"80A6A00F";
    when 16#1F60# => romdata <= X"80A6A000";
    when 16#1F61# => romdata <= X"0280000A";
    when 16#1F62# => romdata <= X"8606BFFF";
    when 16#1F63# => romdata <= X"8406001A";
    when 16#1F64# => romdata <= X"82007FFF";
    when 16#1F65# => romdata <= X"C8084000";
    when 16#1F66# => romdata <= X"8400BFFF";
    when 16#1F67# => romdata <= X"8600FFFF";
    when 16#1F68# => romdata <= X"80A0FFFF";
    when 16#1F69# => romdata <= X"12BFFFFB";
    when 16#1F6A# => romdata <= X"C8288000";
    when 16#1F6B# => romdata <= X"81C7E008";
    when 16#1F6C# => romdata <= X"81E80000";
    when 16#1F6D# => romdata <= X"80A6A00F";
    when 16#1F6E# => romdata <= X"1880000D";
    when 16#1F6F# => romdata <= X"82164018";
    when 16#1F70# => romdata <= X"80A0E000";
    when 16#1F71# => romdata <= X"02BFFFFA";
    when 16#1F72# => romdata <= X"82102000";
    when 16#1F73# => romdata <= X"C4090001";
    when 16#1F74# => romdata <= X"C42B4001";
    when 16#1F75# => romdata <= X"82006001";
    when 16#1F76# => romdata <= X"80A04003";
    when 16#1F77# => romdata <= X"32BFFFFD";
    when 16#1F78# => romdata <= X"C4090001";
    when 16#1F79# => romdata <= X"81C7E008";
    when 16#1F7A# => romdata <= X"81E80000";
    when 16#1F7B# => romdata <= X"80886003";
    when 16#1F7C# => romdata <= X"12BFFFF5";
    when 16#1F7D# => romdata <= X"80A0E000";
    when 16#1F7E# => romdata <= X"8610001A";
    when 16#1F7F# => romdata <= X"84100019";
    when 16#1F80# => romdata <= X"82100018";
    when 16#1F81# => romdata <= X"C8008000";
    when 16#1F82# => romdata <= X"C8204000";
    when 16#1F83# => romdata <= X"8600FFF0";
    when 16#1F84# => romdata <= X"80A0E00F";
    when 16#1F85# => romdata <= X"C800A004";
    when 16#1F86# => romdata <= X"C8206004";
    when 16#1F87# => romdata <= X"C800A008";
    when 16#1F88# => romdata <= X"C8206008";
    when 16#1F89# => romdata <= X"C800A00C";
    when 16#1F8A# => romdata <= X"C820600C";
    when 16#1F8B# => romdata <= X"8400A010";
    when 16#1F8C# => romdata <= X"18BFFFF5";
    when 16#1F8D# => romdata <= X"82006010";
    when 16#1F8E# => romdata <= X"B406BFF0";
    when 16#1F8F# => romdata <= X"9B36A004";
    when 16#1F90# => romdata <= X"832B6004";
    when 16#1F91# => romdata <= X"9A036001";
    when 16#1F92# => romdata <= X"B4268001";
    when 16#1F93# => romdata <= X"9B2B6004";
    when 16#1F94# => romdata <= X"80A6A003";
    when 16#1F95# => romdata <= X"8806400D";
    when 16#1F96# => romdata <= X"8610001A";
    when 16#1F97# => romdata <= X"08BFFFD9";
    when 16#1F98# => romdata <= X"9A06000D";
    when 16#1F99# => romdata <= X"82102000";
    when 16#1F9A# => romdata <= X"C4010001";
    when 16#1F9B# => romdata <= X"C4234001";
    when 16#1F9C# => romdata <= X"82006004";
    when 16#1F9D# => romdata <= X"84268001";
    when 16#1F9E# => romdata <= X"80A0A003";
    when 16#1F9F# => romdata <= X"38BFFFFC";
    when 16#1FA0# => romdata <= X"C4010001";
    when 16#1FA1# => romdata <= X"B406BFFC";
    when 16#1FA2# => romdata <= X"8336A002";
    when 16#1FA3# => romdata <= X"87286002";
    when 16#1FA4# => romdata <= X"82006001";
    when 16#1FA5# => romdata <= X"86268003";
    when 16#1FA6# => romdata <= X"83286002";
    when 16#1FA7# => romdata <= X"88010001";
    when 16#1FA8# => romdata <= X"10BFFFC8";
    when 16#1FA9# => romdata <= X"9A034001";
    when 16#1FAA# => romdata <= X"9DE3BFA0";
    when 16#1FAB# => romdata <= X"860E60FF";
    when 16#1FAC# => romdata <= X"80A6A003";
    when 16#1FAD# => romdata <= X"0880002A";
    when 16#1FAE# => romdata <= X"84100018";
    when 16#1FAF# => romdata <= X"808E2003";
    when 16#1FB0# => romdata <= X"3280002A";
    when 16#1FB1# => romdata <= X"82102000";
    when 16#1FB2# => romdata <= X"8328E008";
    when 16#1FB3# => romdata <= X"82104003";
    when 16#1FB4# => romdata <= X"80A6A00F";
    when 16#1FB5# => romdata <= X"85286010";
    when 16#1FB6# => romdata <= X"9A100018";
    when 16#1FB7# => romdata <= X"84108001";
    when 16#1FB8# => romdata <= X"8810001A";
    when 16#1FB9# => romdata <= X"08800011";
    when 16#1FBA# => romdata <= X"82100018";
    when 16#1FBB# => romdata <= X"C4204000";
    when 16#1FBC# => romdata <= X"C4206004";
    when 16#1FBD# => romdata <= X"C4206008";
    when 16#1FBE# => romdata <= X"C420600C";
    when 16#1FBF# => romdata <= X"88013FF0";
    when 16#1FC0# => romdata <= X"80A1200F";
    when 16#1FC1# => romdata <= X"18BFFFFA";
    when 16#1FC2# => romdata <= X"82006010";
    when 16#1FC3# => romdata <= X"8206BFF0";
    when 16#1FC4# => romdata <= X"B408600F";
    when 16#1FC5# => romdata <= X"9A087FF0";
    when 16#1FC6# => romdata <= X"80A6A003";
    when 16#1FC7# => romdata <= X"9A036010";
    when 16#1FC8# => romdata <= X"0880000E";
    when 16#1FC9# => romdata <= X"9A06000D";
    when 16#1FCA# => romdata <= X"82102000";
    when 16#1FCB# => romdata <= X"C4234001";
    when 16#1FCC# => romdata <= X"82006004";
    when 16#1FCD# => romdata <= X"88268001";
    when 16#1FCE# => romdata <= X"80A12003";
    when 16#1FCF# => romdata <= X"38BFFFFD";
    when 16#1FD0# => romdata <= X"C4234001";
    when 16#1FD1# => romdata <= X"8206BFFC";
    when 16#1FD2# => romdata <= X"B4086003";
    when 16#1FD3# => romdata <= X"82087FFC";
    when 16#1FD4# => romdata <= X"82006004";
    when 16#1FD5# => romdata <= X"9A034001";
    when 16#1FD6# => romdata <= X"8410000D";
    when 16#1FD7# => romdata <= X"80A6A000";
    when 16#1FD8# => romdata <= X"02800007";
    when 16#1FD9# => romdata <= X"82102000";
    when 16#1FDA# => romdata <= X"C6288001";
    when 16#1FDB# => romdata <= X"82006001";
    when 16#1FDC# => romdata <= X"80A0401A";
    when 16#1FDD# => romdata <= X"32BFFFFE";
    when 16#1FDE# => romdata <= X"C6288001";
    when 16#1FDF# => romdata <= X"81C7E008";
    when 16#1FE0# => romdata <= X"81E80000";
    when 16#1FE1# => romdata <= X"80A26000";
    when 16#1FE2# => romdata <= X"02800008";
    when 16#1FE3# => romdata <= X"01000000";
    when 16#1FE4# => romdata <= X"C402204C";
    when 16#1FE5# => romdata <= X"C2026004";
    when 16#1FE6# => romdata <= X"83286002";
    when 16#1FE7# => romdata <= X"C6008001";
    when 16#1FE8# => romdata <= X"C6224000";
    when 16#1FE9# => romdata <= X"D2208001";
    when 16#1FEA# => romdata <= X"81C3E008";
    when 16#1FEB# => romdata <= X"01000000";
    when 16#1FEC# => romdata <= X"82100008";
    when 16#1FED# => romdata <= X"053FFFC0";
    when 16#1FEE# => romdata <= X"808A0002";
    when 16#1FEF# => romdata <= X"12800004";
    when 16#1FF0# => romdata <= X"90102000";
    when 16#1FF1# => romdata <= X"83286010";
    when 16#1FF2# => romdata <= X"90102010";
    when 16#1FF3# => romdata <= X"053FC000";
    when 16#1FF4# => romdata <= X"80884002";
    when 16#1FF5# => romdata <= X"12800004";
    when 16#1FF6# => romdata <= X"053C0000";
    when 16#1FF7# => romdata <= X"90022008";
    when 16#1FF8# => romdata <= X"83286008";
    when 16#1FF9# => romdata <= X"80884002";
    when 16#1FFA# => romdata <= X"12800004";
    when 16#1FFB# => romdata <= X"05300000";
    when 16#1FFC# => romdata <= X"90022004";
    when 16#1FFD# => romdata <= X"83286004";
    when 16#1FFE# => romdata <= X"80884002";
    when 16#1FFF# => romdata <= X"12800005";
    when 16#2000# => romdata <= X"80A06000";
    when 16#2001# => romdata <= X"90022002";
    when 16#2002# => romdata <= X"83286002";
    when 16#2003# => romdata <= X"80A06000";
    when 16#2004# => romdata <= X"06800005";
    when 16#2005# => romdata <= X"05100000";
    when 16#2006# => romdata <= X"80884002";
    when 16#2007# => romdata <= X"02800004";
    when 16#2008# => romdata <= X"90022001";
    when 16#2009# => romdata <= X"81C3E008";
    when 16#200A# => romdata <= X"01000000";
    when 16#200B# => romdata <= X"81C3E008";
    when 16#200C# => romdata <= X"90102020";
    when 16#200D# => romdata <= X"C2020000";
    when 16#200E# => romdata <= X"80886007";
    when 16#200F# => romdata <= X"0280000C";
    when 16#2010# => romdata <= X"0500003F";
    when 16#2011# => romdata <= X"80886001";
    when 16#2012# => romdata <= X"12800007";
    when 16#2013# => romdata <= X"84102000";
    when 16#2014# => romdata <= X"80886002";
    when 16#2015# => romdata <= X"1280002C";
    when 16#2016# => romdata <= X"84102002";
    when 16#2017# => romdata <= X"83306002";
    when 16#2018# => romdata <= X"C2220000";
    when 16#2019# => romdata <= X"81C3E008";
    when 16#201A# => romdata <= X"90100002";
    when 16#201B# => romdata <= X"8410A3FF";
    when 16#201C# => romdata <= X"80884002";
    when 16#201D# => romdata <= X"0280001B";
    when 16#201E# => romdata <= X"84102000";
    when 16#201F# => romdata <= X"808860FF";
    when 16#2020# => romdata <= X"12800005";
    when 16#2021# => romdata <= X"8088600F";
    when 16#2022# => romdata <= X"8400A008";
    when 16#2023# => romdata <= X"83306008";
    when 16#2024# => romdata <= X"8088600F";
    when 16#2025# => romdata <= X"12800005";
    when 16#2026# => romdata <= X"80886003";
    when 16#2027# => romdata <= X"8400A004";
    when 16#2028# => romdata <= X"83306004";
    when 16#2029# => romdata <= X"80886003";
    when 16#202A# => romdata <= X"12800005";
    when 16#202B# => romdata <= X"80886001";
    when 16#202C# => romdata <= X"8400A002";
    when 16#202D# => romdata <= X"83306002";
    when 16#202E# => romdata <= X"80886001";
    when 16#202F# => romdata <= X"32800007";
    when 16#2030# => romdata <= X"C2220000";
    when 16#2031# => romdata <= X"83306001";
    when 16#2032# => romdata <= X"80A06000";
    when 16#2033# => romdata <= X"0280000B";
    when 16#2034# => romdata <= X"8400A001";
    when 16#2035# => romdata <= X"C2220000";
    when 16#2036# => romdata <= X"81C3E008";
    when 16#2037# => romdata <= X"90100002";
    when 16#2038# => romdata <= X"83306010";
    when 16#2039# => romdata <= X"808860FF";
    when 16#203A# => romdata <= X"12BFFFEA";
    when 16#203B# => romdata <= X"84102010";
    when 16#203C# => romdata <= X"10BFFFE7";
    when 16#203D# => romdata <= X"8400A008";
    when 16#203E# => romdata <= X"84102020";
    when 16#203F# => romdata <= X"81C3E008";
    when 16#2040# => romdata <= X"90100002";
    when 16#2041# => romdata <= X"83306001";
    when 16#2042# => romdata <= X"84102001";
    when 16#2043# => romdata <= X"C2220000";
    when 16#2044# => romdata <= X"81C3E008";
    when 16#2045# => romdata <= X"90100002";
    when 16#2046# => romdata <= X"9DE3BFA0";
    when 16#2047# => romdata <= X"82100018";
    when 16#2048# => romdata <= X"C4066010";
    when 16#2049# => romdata <= X"F0062010";
    when 16#204A# => romdata <= X"B0A60002";
    when 16#204B# => romdata <= X"12800011";
    when 16#204C# => romdata <= X"8400A004";
    when 16#204D# => romdata <= X"8528A002";
    when 16#204E# => romdata <= X"86064002";
    when 16#204F# => romdata <= X"84004002";
    when 16#2050# => romdata <= X"8600E004";
    when 16#2051# => romdata <= X"8400A004";
    when 16#2052# => romdata <= X"82006014";
    when 16#2053# => romdata <= X"8400BFFC";
    when 16#2054# => romdata <= X"8600FFFC";
    when 16#2055# => romdata <= X"DA008000";
    when 16#2056# => romdata <= X"C800C000";
    when 16#2057# => romdata <= X"80A34004";
    when 16#2058# => romdata <= X"12800006";
    when 16#2059# => romdata <= X"80A04002";
    when 16#205A# => romdata <= X"0ABFFFFA";
    when 16#205B# => romdata <= X"8400BFFC";
    when 16#205C# => romdata <= X"81C7E008";
    when 16#205D# => romdata <= X"81E80000";
    when 16#205E# => romdata <= X"80A34004";
    when 16#205F# => romdata <= X"B0602000";
    when 16#2060# => romdata <= X"B0162001";
    when 16#2061# => romdata <= X"81C7E008";
    when 16#2062# => romdata <= X"81E80000";
    when 16#2063# => romdata <= X"031FFC00";
    when 16#2064# => romdata <= X"053F3000";
    when 16#2065# => romdata <= X"820A0001";
    when 16#2066# => romdata <= X"82004002";
    when 16#2067# => romdata <= X"80A06000";
    when 16#2068# => romdata <= X"04800008";
    when 16#2069# => romdata <= X"9C03BF98";
    when 16#206A# => romdata <= X"84100001";
    when 16#206B# => romdata <= X"86102000";
    when 16#206C# => romdata <= X"C43BA060";
    when 16#206D# => romdata <= X"C11BA060";
    when 16#206E# => romdata <= X"81C3E008";
    when 16#206F# => romdata <= X"9C23BF98";
    when 16#2070# => romdata <= X"82200001";
    when 16#2071# => romdata <= X"83386014";
    when 16#2072# => romdata <= X"80A06013";
    when 16#2073# => romdata <= X"04800011";
    when 16#2074# => romdata <= X"09000200";
    when 16#2075# => romdata <= X"82007FEC";
    when 16#2076# => romdata <= X"80A0601E";
    when 16#2077# => romdata <= X"04800008";
    when 16#2078# => romdata <= X"88102001";
    when 16#2079# => romdata <= X"84102000";
    when 16#207A# => romdata <= X"86100004";
    when 16#207B# => romdata <= X"C43BA060";
    when 16#207C# => romdata <= X"C11BA060";
    when 16#207D# => romdata <= X"81C3E008";
    when 16#207E# => romdata <= X"9C23BF98";
    when 16#207F# => romdata <= X"82380001";
    when 16#2080# => romdata <= X"84102000";
    when 16#2081# => romdata <= X"89290001";
    when 16#2082# => romdata <= X"10BFFFF9";
    when 16#2083# => romdata <= X"86100004";
    when 16#2084# => romdata <= X"86102000";
    when 16#2085# => romdata <= X"85390001";
    when 16#2086# => romdata <= X"C43BA060";
    when 16#2087# => romdata <= X"C11BA060";
    when 16#2088# => romdata <= X"81C3E008";
    when 16#2089# => romdata <= X"9C23BF98";
    when 16#208A# => romdata <= X"9DE3BF98";
    when 16#208B# => romdata <= X"E0062010";
    when 16#208C# => romdata <= X"A0042004";
    when 16#208D# => romdata <= X"A12C2002";
    when 16#208E# => romdata <= X"E2060010";
    when 16#208F# => romdata <= X"7FFFFF5D";
    when 16#2090# => romdata <= X"90100011";
    when 16#2091# => romdata <= X"82102020";
    when 16#2092# => romdata <= X"82204008";
    when 16#2093# => romdata <= X"C2264000";
    when 16#2094# => romdata <= X"A0060010";
    when 16#2095# => romdata <= X"80A2200A";
    when 16#2096# => romdata <= X"14800013";
    when 16#2097# => romdata <= X"B0062014";
    when 16#2098# => romdata <= X"8410200B";
    when 16#2099# => romdata <= X"80A60010";
    when 16#209A# => romdata <= X"84208008";
    when 16#209B# => romdata <= X"1A800004";
    when 16#209C# => romdata <= X"82102000";
    when 16#209D# => romdata <= X"C2043FFC";
    when 16#209E# => romdata <= X"83304002";
    when 16#209F# => romdata <= X"9B344002";
    when 16#20A0# => romdata <= X"90022015";
    when 16#20A1# => romdata <= X"090FFC00";
    when 16#20A2# => romdata <= X"A32C4008";
    when 16#20A3# => romdata <= X"84134004";
    when 16#20A4# => romdata <= X"86104011";
    when 16#20A5# => romdata <= X"C43FBFF8";
    when 16#20A6# => romdata <= X"C11FBFF8";
    when 16#20A7# => romdata <= X"81C7E008";
    when 16#20A8# => romdata <= X"81E80000";
    when 16#20A9# => romdata <= X"80A60010";
    when 16#20AA# => romdata <= X"0A80001E";
    when 16#20AB# => romdata <= X"82102000";
    when 16#20AC# => romdata <= X"90823FF5";
    when 16#20AD# => romdata <= X"02800015";
    when 16#20AE# => romdata <= X"090FFC00";
    when 16#20AF# => romdata <= X"84102020";
    when 16#20B0# => romdata <= X"80A40018";
    when 16#20B1# => romdata <= X"84208008";
    when 16#20B2# => romdata <= X"08800004";
    when 16#20B3# => romdata <= X"88102000";
    when 16#20B4# => romdata <= X"C8043FFC";
    when 16#20B5# => romdata <= X"89310002";
    when 16#20B6# => romdata <= X"9B284008";
    when 16#20B7# => romdata <= X"83304002";
    when 16#20B8# => romdata <= X"050FFC00";
    when 16#20B9# => romdata <= X"912C4008";
    when 16#20BA# => romdata <= X"8611000D";
    when 16#20BB# => romdata <= X"90120002";
    when 16#20BC# => romdata <= X"84120001";
    when 16#20BD# => romdata <= X"C43FBFF8";
    when 16#20BE# => romdata <= X"C11FBFF8";
    when 16#20BF# => romdata <= X"81C7E008";
    when 16#20C0# => romdata <= X"81E80000";
    when 16#20C1# => romdata <= X"090FFC00";
    when 16#20C2# => romdata <= X"86100001";
    when 16#20C3# => romdata <= X"84144004";
    when 16#20C4# => romdata <= X"C43FBFF8";
    when 16#20C5# => romdata <= X"C11FBFF8";
    when 16#20C6# => romdata <= X"81C7E008";
    when 16#20C7# => romdata <= X"81E80000";
    when 16#20C8# => romdata <= X"C2043FFC";
    when 16#20C9# => romdata <= X"90823FF5";
    when 16#20CA# => romdata <= X"02BFFFF7";
    when 16#20CB# => romdata <= X"A0043FFC";
    when 16#20CC# => romdata <= X"10BFFFE4";
    when 16#20CD# => romdata <= X"84102020";
    when 16#20CE# => romdata <= X"9DE3BF88";
    when 16#20CF# => romdata <= X"9207BFFC";
    when 16#20D0# => romdata <= X"7FFFFFBA";
    when 16#20D1# => romdata <= X"90100018";
    when 16#20D2# => romdata <= X"91A00020";
    when 16#20D3# => romdata <= X"9207BFF8";
    when 16#20D4# => romdata <= X"90100019";
    when 16#20D5# => romdata <= X"C327BFF0";
    when 16#20D6# => romdata <= X"7FFFFFB4";
    when 16#20D7# => romdata <= X"D127BFF4";
    when 16#20D8# => romdata <= X"C6062010";
    when 16#20D9# => romdata <= X"C4066010";
    when 16#20DA# => romdata <= X"C207BFF8";
    when 16#20DB# => romdata <= X"C807BFFC";
    when 16#20DC# => romdata <= X"82210001";
    when 16#20DD# => romdata <= X"8420C002";
    when 16#20DE# => romdata <= X"D107BFF4";
    when 16#20DF# => romdata <= X"8528A005";
    when 16#20E0# => romdata <= X"D307BFF0";
    when 16#20E1# => romdata <= X"82004002";
    when 16#20E2# => romdata <= X"80A06000";
    when 16#20E3# => romdata <= X"0480000C";
    when 16#20E4# => romdata <= X"99A00020";
    when 16#20E5# => romdata <= X"D127BFEC";
    when 16#20E6# => romdata <= X"83286014";
    when 16#20E7# => romdata <= X"C407BFEC";
    when 16#20E8# => romdata <= X"82004002";
    when 16#20E9# => romdata <= X"C227BFEC";
    when 16#20EA# => romdata <= X"D507BFEC";
    when 16#20EB# => romdata <= X"91A0002A";
    when 16#20EC# => romdata <= X"81A209C0";
    when 16#20ED# => romdata <= X"81C7E008";
    when 16#20EE# => romdata <= X"81E80000";
    when 16#20EF# => romdata <= X"D927BFEC";
    when 16#20F0# => romdata <= X"83286014";
    when 16#20F1# => romdata <= X"C407BFEC";
    when 16#20F2# => romdata <= X"82208001";
    when 16#20F3# => romdata <= X"C227BFEC";
    when 16#20F4# => romdata <= X"D907BFEC";
    when 16#20F5# => romdata <= X"81A0002C";
    when 16#20F6# => romdata <= X"81A209C0";
    when 16#20F7# => romdata <= X"81C7E008";
    when 16#20F8# => romdata <= X"81E80000";
    when 16#20F9# => romdata <= X"80A22017";
    when 16#20FA# => romdata <= X"0480000A";
    when 16#20FB# => romdata <= X"03100032";
    when 16#20FC# => romdata <= X"C11860E0";
    when 16#20FD# => romdata <= X"03100032";
    when 16#20FE# => romdata <= X"D11860E8";
    when 16#20FF# => romdata <= X"90823FFF";
    when 16#2100# => romdata <= X"12BFFFFF";
    when 16#2101# => romdata <= X"81A00948";
    when 16#2102# => romdata <= X"81C3E008";
    when 16#2103# => romdata <= X"01000000";
    when 16#2104# => romdata <= X"912A2003";
    when 16#2105# => romdata <= X"03100032";
    when 16#2106# => romdata <= X"82106150";
    when 16#2107# => romdata <= X"81C3E008";
    when 16#2108# => romdata <= X"C1184008";
    when 16#2109# => romdata <= X"9DE3BFA0";
    when 16#210A# => romdata <= X"C206204C";
    when 16#210B# => romdata <= X"80A06000";
    when 16#210C# => romdata <= X"0280000D";
    when 16#210D# => romdata <= X"A0100018";
    when 16#210E# => romdata <= X"852E6002";
    when 16#210F# => romdata <= X"F0004002";
    when 16#2110# => romdata <= X"80A62000";
    when 16#2111# => romdata <= X"02800013";
    when 16#2112# => romdata <= X"90100010";
    when 16#2113# => romdata <= X"C6060000";
    when 16#2114# => romdata <= X"C6204002";
    when 16#2115# => romdata <= X"C0262010";
    when 16#2116# => romdata <= X"C026200C";
    when 16#2117# => romdata <= X"81C7E008";
    when 16#2118# => romdata <= X"81E80000";
    when 16#2119# => romdata <= X"90100018";
    when 16#211A# => romdata <= X"92102004";
    when 16#211B# => romdata <= X"400004A3";
    when 16#211C# => romdata <= X"94102010";
    when 16#211D# => romdata <= X"D024204C";
    when 16#211E# => romdata <= X"82100008";
    when 16#211F# => romdata <= X"80A22000";
    when 16#2120# => romdata <= X"12BFFFEE";
    when 16#2121# => romdata <= X"B0102000";
    when 16#2122# => romdata <= X"81C7E008";
    when 16#2123# => romdata <= X"81E80000";
    when 16#2124# => romdata <= X"92102001";
    when 16#2125# => romdata <= X"A0102001";
    when 16#2126# => romdata <= X"A12C0019";
    when 16#2127# => romdata <= X"94042005";
    when 16#2128# => romdata <= X"40000496";
    when 16#2129# => romdata <= X"952AA002";
    when 16#212A# => romdata <= X"B0922000";
    when 16#212B# => romdata <= X"02BFFFF7";
    when 16#212C# => romdata <= X"01000000";
    when 16#212D# => romdata <= X"F2262004";
    when 16#212E# => romdata <= X"E0262008";
    when 16#212F# => romdata <= X"C0262010";
    when 16#2130# => romdata <= X"C026200C";
    when 16#2131# => romdata <= X"81C7E008";
    when 16#2132# => romdata <= X"81E80000";
    when 16#2133# => romdata <= X"9DE3BF90";
    when 16#2134# => romdata <= X"92102001";
    when 16#2135# => romdata <= X"90100018";
    when 16#2136# => romdata <= X"F227BFF0";
    when 16#2137# => romdata <= X"7FFFFFD2";
    when 16#2138# => romdata <= X"F427BFF4";
    when 16#2139# => romdata <= X"053FFC00";
    when 16#213A# => romdata <= X"842E4002";
    when 16#213B# => romdata <= X"C427BFF8";
    when 16#213C# => romdata <= X"07200000";
    when 16#213D# => romdata <= X"A210001A";
    when 16#213E# => romdata <= X"822E4003";
    when 16#213F# => romdata <= X"A5306014";
    when 16#2140# => romdata <= X"80A4A000";
    when 16#2141# => romdata <= X"02800005";
    when 16#2142# => romdata <= X"B0100008";
    when 16#2143# => romdata <= X"07000400";
    when 16#2144# => romdata <= X"84108003";
    when 16#2145# => romdata <= X"C427BFF8";
    when 16#2146# => romdata <= X"80A46000";
    when 16#2147# => romdata <= X"0280001E";
    when 16#2148# => romdata <= X"01000000";
    when 16#2149# => romdata <= X"E227BFFC";
    when 16#214A# => romdata <= X"7FFFFEC3";
    when 16#214B# => romdata <= X"9007BFFC";
    when 16#214C# => romdata <= X"80A22000";
    when 16#214D# => romdata <= X"1280002A";
    when 16#214E# => romdata <= X"C207BFF8";
    when 16#214F# => romdata <= X"C207BFFC";
    when 16#2150# => romdata <= X"C2262014";
    when 16#2151# => romdata <= X"C207BFF8";
    when 16#2152# => romdata <= X"80A00001";
    when 16#2153# => romdata <= X"C2262018";
    when 16#2154# => romdata <= X"A0402000";
    when 16#2155# => romdata <= X"A0042001";
    when 16#2156# => romdata <= X"80A4A000";
    when 16#2157# => romdata <= X"12800018";
    when 16#2158# => romdata <= X"E0262010";
    when 16#2159# => romdata <= X"90023BCE";
    when 16#215A# => romdata <= X"82042003";
    when 16#215B# => romdata <= X"D026C000";
    when 16#215C# => romdata <= X"83286002";
    when 16#215D# => romdata <= X"82060001";
    when 16#215E# => romdata <= X"7FFFFE8E";
    when 16#215F# => romdata <= X"D0006004";
    when 16#2160# => romdata <= X"A12C2005";
    when 16#2161# => romdata <= X"A0240008";
    when 16#2162# => romdata <= X"E0270000";
    when 16#2163# => romdata <= X"81C7E008";
    when 16#2164# => romdata <= X"81E80000";
    when 16#2165# => romdata <= X"7FFFFEA8";
    when 16#2166# => romdata <= X"9007BFF8";
    when 16#2167# => romdata <= X"C207BFF8";
    when 16#2168# => romdata <= X"C2262014";
    when 16#2169# => romdata <= X"82102001";
    when 16#216A# => romdata <= X"C2262010";
    when 16#216B# => romdata <= X"90022020";
    when 16#216C# => romdata <= X"80A4A000";
    when 16#216D# => romdata <= X"02BFFFEC";
    when 16#216E# => romdata <= X"A0102001";
    when 16#216F# => romdata <= X"A404BBCD";
    when 16#2170# => romdata <= X"A4048008";
    when 16#2171# => romdata <= X"E426C000";
    when 16#2172# => romdata <= X"82102035";
    when 16#2173# => romdata <= X"90204008";
    when 16#2174# => romdata <= X"D0270000";
    when 16#2175# => romdata <= X"81C7E008";
    when 16#2176# => romdata <= X"81E80000";
    when 16#2177# => romdata <= X"C607BFFC";
    when 16#2178# => romdata <= X"84200008";
    when 16#2179# => romdata <= X"85284002";
    when 16#217A# => romdata <= X"84108003";
    when 16#217B# => romdata <= X"C4262014";
    when 16#217C# => romdata <= X"83304008";
    when 16#217D# => romdata <= X"10BFFFD5";
    when 16#217E# => romdata <= X"C227BFF8";
    when 16#217F# => romdata <= X"9DE3BFA0";
    when 16#2180# => romdata <= X"E2066010";
    when 16#2181# => romdata <= X"C206A010";
    when 16#2182# => romdata <= X"A2A44001";
    when 16#2183# => romdata <= X"0280004A";
    when 16#2184# => romdata <= X"90100018";
    when 16#2185# => romdata <= X"80A46000";
    when 16#2186# => romdata <= X"06800061";
    when 16#2187# => romdata <= X"82100019";
    when 16#2188# => romdata <= X"A2102000";
    when 16#2189# => romdata <= X"A0066014";
    when 16#218A# => romdata <= X"7FFFFF7F";
    when 16#218B# => romdata <= X"D2066004";
    when 16#218C# => romdata <= X"C8066010";
    when 16#218D# => romdata <= X"D206A010";
    when 16#218E# => romdata <= X"82012004";
    when 16#218F# => romdata <= X"E222200C";
    when 16#2190# => romdata <= X"83286002";
    when 16#2191# => romdata <= X"92026004";
    when 16#2192# => romdata <= X"B2064001";
    when 16#2193# => romdata <= X"932A6002";
    when 16#2194# => romdata <= X"1900003F";
    when 16#2195# => romdata <= X"92068009";
    when 16#2196# => romdata <= X"B2066004";
    when 16#2197# => romdata <= X"92026004";
    when 16#2198# => romdata <= X"981323FF";
    when 16#2199# => romdata <= X"B406A014";
    when 16#219A# => romdata <= X"82022014";
    when 16#219B# => romdata <= X"84102000";
    when 16#219C# => romdata <= X"DA068000";
    when 16#219D# => romdata <= X"C6040000";
    when 16#219E# => romdata <= X"97336010";
    when 16#219F# => romdata <= X"9A0B400C";
    when 16#21A0# => romdata <= X"9530E010";
    when 16#21A1# => romdata <= X"8608C00C";
    when 16#21A2# => romdata <= X"9622800B";
    when 16#21A3# => romdata <= X"8620C00D";
    when 16#21A4# => romdata <= X"8600C002";
    when 16#21A5# => romdata <= X"9B38E010";
    when 16#21A6# => romdata <= X"8402C00D";
    when 16#21A7# => romdata <= X"C6306002";
    when 16#21A8# => romdata <= X"B406A004";
    when 16#21A9# => romdata <= X"C4304000";
    when 16#21AA# => romdata <= X"A0042004";
    when 16#21AB# => romdata <= X"82006004";
    when 16#21AC# => romdata <= X"80A2401A";
    when 16#21AD# => romdata <= X"18BFFFEF";
    when 16#21AE# => romdata <= X"8538A010";
    when 16#21AF# => romdata <= X"80A40019";
    when 16#21B0# => romdata <= X"3A800012";
    when 16#21B1# => romdata <= X"C4007FFC";
    when 16#21B2# => romdata <= X"1900003F";
    when 16#21B3# => romdata <= X"981323FF";
    when 16#21B4# => romdata <= X"C6040000";
    when 16#21B5# => romdata <= X"9B30E010";
    when 16#21B6# => romdata <= X"8608C00C";
    when 16#21B7# => romdata <= X"86008003";
    when 16#21B8# => romdata <= X"8538E010";
    when 16#21B9# => romdata <= X"8400800D";
    when 16#21BA# => romdata <= X"C6306002";
    when 16#21BB# => romdata <= X"A0042004";
    when 16#21BC# => romdata <= X"C4304000";
    when 16#21BD# => romdata <= X"80A64010";
    when 16#21BE# => romdata <= X"82006004";
    when 16#21BF# => romdata <= X"18BFFFF5";
    when 16#21C0# => romdata <= X"8538A010";
    when 16#21C1# => romdata <= X"C4007FFC";
    when 16#21C2# => romdata <= X"80A0A000";
    when 16#21C3# => romdata <= X"12800007";
    when 16#21C4# => romdata <= X"82007FFC";
    when 16#21C5# => romdata <= X"82007FFC";
    when 16#21C6# => romdata <= X"C4004000";
    when 16#21C7# => romdata <= X"80A0A000";
    when 16#21C8# => romdata <= X"02BFFFFD";
    when 16#21C9# => romdata <= X"88013FFF";
    when 16#21CA# => romdata <= X"C8222010";
    when 16#21CB# => romdata <= X"81C7E008";
    when 16#21CC# => romdata <= X"91E80008";
    when 16#21CD# => romdata <= X"82006004";
    when 16#21CE# => romdata <= X"A0066014";
    when 16#21CF# => romdata <= X"83286002";
    when 16#21D0# => romdata <= X"84068001";
    when 16#21D1# => romdata <= X"82064001";
    when 16#21D2# => romdata <= X"8400A004";
    when 16#21D3# => romdata <= X"82006004";
    when 16#21D4# => romdata <= X"82007FFC";
    when 16#21D5# => romdata <= X"8400BFFC";
    when 16#21D6# => romdata <= X"C8004000";
    when 16#21D7# => romdata <= X"C6008000";
    when 16#21D8# => romdata <= X"80A10003";
    when 16#21D9# => romdata <= X"1280000B";
    when 16#21DA# => romdata <= X"80A40001";
    when 16#21DB# => romdata <= X"0ABFFFFA";
    when 16#21DC# => romdata <= X"82007FFC";
    when 16#21DD# => romdata <= X"7FFFFF2C";
    when 16#21DE# => romdata <= X"92102000";
    when 16#21DF# => romdata <= X"82102001";
    when 16#21E0# => romdata <= X"C0222014";
    when 16#21E1# => romdata <= X"C2222010";
    when 16#21E2# => romdata <= X"81C7E008";
    when 16#21E3# => romdata <= X"91E80008";
    when 16#21E4# => romdata <= X"80A10003";
    when 16#21E5# => romdata <= X"1ABFFFA5";
    when 16#21E6# => romdata <= X"82100019";
    when 16#21E7# => romdata <= X"A2102001";
    when 16#21E8# => romdata <= X"B210001A";
    when 16#21E9# => romdata <= X"B4100001";
    when 16#21EA# => romdata <= X"10BFFFA0";
    when 16#21EB# => romdata <= X"A0066014";
    when 16#21EC# => romdata <= X"9DE3BFA0";
    when 16#21ED# => romdata <= X"E0066010";
    when 16#21EE# => romdata <= X"C2066008";
    when 16#21EF# => romdata <= X"A0042001";
    when 16#21F0# => romdata <= X"A33EA005";
    when 16#21F1# => romdata <= X"A4100018";
    when 16#21F2# => romdata <= X"A0040011";
    when 16#21F3# => romdata <= X"80A40001";
    when 16#21F4# => romdata <= X"04800006";
    when 16#21F5# => romdata <= X"D2066004";
    when 16#21F6# => romdata <= X"83286001";
    when 16#21F7# => romdata <= X"80A40001";
    when 16#21F8# => romdata <= X"14BFFFFE";
    when 16#21F9# => romdata <= X"92026001";
    when 16#21FA# => romdata <= X"7FFFFF0F";
    when 16#21FB# => romdata <= X"90100012";
    when 16#21FC# => romdata <= X"80A46000";
    when 16#21FD# => romdata <= X"0480000C";
    when 16#21FE# => romdata <= X"82022014";
    when 16#21FF# => romdata <= X"84102000";
    when 16#2200# => romdata <= X"C0204000";
    when 16#2201# => romdata <= X"8400A001";
    when 16#2202# => romdata <= X"80A08011";
    when 16#2203# => romdata <= X"12BFFFFD";
    when 16#2204# => romdata <= X"82006004";
    when 16#2205# => romdata <= X"8200A004";
    when 16#2206# => romdata <= X"83286002";
    when 16#2207# => romdata <= X"82020001";
    when 16#2208# => romdata <= X"82006004";
    when 16#2209# => romdata <= X"C8066010";
    when 16#220A# => romdata <= X"88012004";
    when 16#220B# => romdata <= X"B48EA01F";
    when 16#220C# => romdata <= X"89292002";
    when 16#220D# => romdata <= X"84066014";
    when 16#220E# => romdata <= X"88064004";
    when 16#220F# => romdata <= X"0280001C";
    when 16#2210# => romdata <= X"88012004";
    when 16#2211# => romdata <= X"98102020";
    when 16#2212# => romdata <= X"86102000";
    when 16#2213# => romdata <= X"9823001A";
    when 16#2214# => romdata <= X"DA008000";
    when 16#2215# => romdata <= X"9B2B401A";
    when 16#2216# => romdata <= X"8610C00D";
    when 16#2217# => romdata <= X"C6204000";
    when 16#2218# => romdata <= X"82006004";
    when 16#2219# => romdata <= X"C6008000";
    when 16#221A# => romdata <= X"8400A004";
    when 16#221B# => romdata <= X"80A10002";
    when 16#221C# => romdata <= X"18BFFFF8";
    when 16#221D# => romdata <= X"8730C00C";
    when 16#221E# => romdata <= X"C6204000";
    when 16#221F# => romdata <= X"80A00003";
    when 16#2220# => romdata <= X"A0400010";
    when 16#2221# => romdata <= X"C404A04C";
    when 16#2222# => romdata <= X"C2066004";
    when 16#2223# => romdata <= X"83286002";
    when 16#2224# => romdata <= X"C6008001";
    when 16#2225# => romdata <= X"C6264000";
    when 16#2226# => romdata <= X"A0043FFF";
    when 16#2227# => romdata <= X"F2208001";
    when 16#2228# => romdata <= X"E0222010";
    when 16#2229# => romdata <= X"81C7E008";
    when 16#222A# => romdata <= X"91E80008";
    when 16#222B# => romdata <= X"C6008000";
    when 16#222C# => romdata <= X"C6204000";
    when 16#222D# => romdata <= X"8400A004";
    when 16#222E# => romdata <= X"80A10002";
    when 16#222F# => romdata <= X"08BFFFF2";
    when 16#2230# => romdata <= X"82006004";
    when 16#2231# => romdata <= X"C6008000";
    when 16#2232# => romdata <= X"C6204000";
    when 16#2233# => romdata <= X"8400A004";
    when 16#2234# => romdata <= X"80A10002";
    when 16#2235# => romdata <= X"18BFFFF6";
    when 16#2236# => romdata <= X"82006004";
    when 16#2237# => romdata <= X"10BFFFEB";
    when 16#2238# => romdata <= X"C404A04C";
    when 16#2239# => romdata <= X"9DE3BF98";
    when 16#223A# => romdata <= X"E0066010";
    when 16#223B# => romdata <= X"E206A010";
    when 16#223C# => romdata <= X"80A40011";
    when 16#223D# => romdata <= X"06800080";
    when 16#223E# => romdata <= X"90100018";
    when 16#223F# => romdata <= X"82100011";
    when 16#2240# => romdata <= X"A2100010";
    when 16#2241# => romdata <= X"A0100001";
    when 16#2242# => romdata <= X"C2066008";
    when 16#2243# => romdata <= X"AC040011";
    when 16#2244# => romdata <= X"80A58001";
    when 16#2245# => romdata <= X"04800003";
    when 16#2246# => romdata <= X"D2066004";
    when 16#2247# => romdata <= X"92026001";
    when 16#2248# => romdata <= X"7FFFFEC1";
    when 16#2249# => romdata <= X"AE05A004";
    when 16#224A# => romdata <= X"B6022014";
    when 16#224B# => romdata <= X"AF2DE002";
    when 16#224C# => romdata <= X"AE020017";
    when 16#224D# => romdata <= X"AE05E004";
    when 16#224E# => romdata <= X"80A6C017";
    when 16#224F# => romdata <= X"1A800008";
    when 16#2250# => romdata <= X"B0100008";
    when 16#2251# => romdata <= X"8210001B";
    when 16#2252# => romdata <= X"C0204000";
    when 16#2253# => romdata <= X"82006004";
    when 16#2254# => romdata <= X"80A5C001";
    when 16#2255# => romdata <= X"38BFFFFE";
    when 16#2256# => romdata <= X"C0204000";
    when 16#2257# => romdata <= X"AA046004";
    when 16#2258# => romdata <= X"AB2D6002";
    when 16#2259# => romdata <= X"AA064015";
    when 16#225A# => romdata <= X"B2066014";
    when 16#225B# => romdata <= X"F227BFF8";
    when 16#225C# => romdata <= X"B8042004";
    when 16#225D# => romdata <= X"BA06A014";
    when 16#225E# => romdata <= X"B92F2002";
    when 16#225F# => romdata <= X"B806801C";
    when 16#2260# => romdata <= X"B8072004";
    when 16#2261# => romdata <= X"80A7401C";
    when 16#2262# => romdata <= X"1A800047";
    when 16#2263# => romdata <= X"AA056004";
    when 16#2264# => romdata <= X"2300003F";
    when 16#2265# => romdata <= X"A21463FF";
    when 16#2266# => romdata <= X"C2074000";
    when 16#2267# => romdata <= X"84884011";
    when 16#2268# => romdata <= X"0280001D";
    when 16#2269# => romdata <= X"C427BFFC";
    when 16#226A# => romdata <= X"F407BFF8";
    when 16#226B# => romdata <= X"A010001B";
    when 16#226C# => romdata <= X"B2102000";
    when 16#226D# => romdata <= X"E8068000";
    when 16#226E# => romdata <= X"D207BFFC";
    when 16#226F# => romdata <= X"4000041F";
    when 16#2270# => romdata <= X"900D0011";
    when 16#2271# => romdata <= X"E6040000";
    when 16#2272# => romdata <= X"D207BFFC";
    when 16#2273# => romdata <= X"A40CC011";
    when 16#2274# => romdata <= X"A4020012";
    when 16#2275# => romdata <= X"40000419";
    when 16#2276# => romdata <= X"91352010";
    when 16#2277# => romdata <= X"A4048019";
    when 16#2278# => romdata <= X"A734E010";
    when 16#2279# => romdata <= X"8334A010";
    when 16#227A# => romdata <= X"A6020013";
    when 16#227B# => romdata <= X"B204C001";
    when 16#227C# => romdata <= X"E4342002";
    when 16#227D# => romdata <= X"B406A004";
    when 16#227E# => romdata <= X"F2340000";
    when 16#227F# => romdata <= X"80A5401A";
    when 16#2280# => romdata <= X"A0042004";
    when 16#2281# => romdata <= X"18BFFFEC";
    when 16#2282# => romdata <= X"B3366010";
    when 16#2283# => romdata <= X"F2240000";
    when 16#2284# => romdata <= X"C2074000";
    when 16#2285# => romdata <= X"83306010";
    when 16#2286# => romdata <= X"80A06000";
    when 16#2287# => romdata <= X"0280001E";
    when 16#2288# => romdata <= X"C227BFFC";
    when 16#2289# => romdata <= X"F206C000";
    when 16#228A# => romdata <= X"F407BFF8";
    when 16#228B# => romdata <= X"A4100019";
    when 16#228C# => romdata <= X"A010001B";
    when 16#228D# => romdata <= X"A6102000";
    when 16#228E# => romdata <= X"E8068000";
    when 16#228F# => romdata <= X"D007BFFC";
    when 16#2290# => romdata <= X"920D0011";
    when 16#2291# => romdata <= X"400003FD";
    when 16#2292# => romdata <= X"A534A010";
    when 16#2293# => romdata <= X"A604C008";
    when 16#2294# => romdata <= X"A604C012";
    when 16#2295# => romdata <= X"F2342002";
    when 16#2296# => romdata <= X"D007BFFC";
    when 16#2297# => romdata <= X"E6340000";
    when 16#2298# => romdata <= X"93352010";
    when 16#2299# => romdata <= X"400003F5";
    when 16#229A# => romdata <= X"A734E010";
    when 16#229B# => romdata <= X"A0042004";
    when 16#229C# => romdata <= X"E4040000";
    when 16#229D# => romdata <= X"B406A004";
    when 16#229E# => romdata <= X"B20C8011";
    when 16#229F# => romdata <= X"80A5401A";
    when 16#22A0# => romdata <= X"B2020019";
    when 16#22A1# => romdata <= X"B2064013";
    when 16#22A2# => romdata <= X"18BFFFEC";
    when 16#22A3# => romdata <= X"A7366010";
    when 16#22A4# => romdata <= X"F2240000";
    when 16#22A5# => romdata <= X"BA076004";
    when 16#22A6# => romdata <= X"80A7001D";
    when 16#22A7# => romdata <= X"18BFFFBF";
    when 16#22A8# => romdata <= X"B606E004";
    when 16#22A9# => romdata <= X"80A5A000";
    when 16#22AA# => romdata <= X"24800011";
    when 16#22AB# => romdata <= X"EC262010";
    when 16#22AC# => romdata <= X"C205FFFC";
    when 16#22AD# => romdata <= X"80A06000";
    when 16#22AE# => romdata <= X"02800009";
    when 16#22AF# => romdata <= X"AE05FFFC";
    when 16#22B0# => romdata <= X"EC262010";
    when 16#22B1# => romdata <= X"81C7E008";
    when 16#22B2# => romdata <= X"81E80000";
    when 16#22B3# => romdata <= X"C205C000";
    when 16#22B4# => romdata <= X"80A06000";
    when 16#22B5# => romdata <= X"32800006";
    when 16#22B6# => romdata <= X"EC262010";
    when 16#22B7# => romdata <= X"AC85BFFF";
    when 16#22B8# => romdata <= X"12BFFFFB";
    when 16#22B9# => romdata <= X"AE05FFFC";
    when 16#22BA# => romdata <= X"EC262010";
    when 16#22BB# => romdata <= X"81C7E008";
    when 16#22BC# => romdata <= X"81E80000";
    when 16#22BD# => romdata <= X"82100019";
    when 16#22BE# => romdata <= X"B210001A";
    when 16#22BF# => romdata <= X"10BFFF83";
    when 16#22C0# => romdata <= X"B4100001";
    when 16#22C1# => romdata <= X"9DE3BFA0";
    when 16#22C2# => romdata <= X"92102001";
    when 16#22C3# => romdata <= X"7FFFFE46";
    when 16#22C4# => romdata <= X"90100018";
    when 16#22C5# => romdata <= X"82102001";
    when 16#22C6# => romdata <= X"F2222014";
    when 16#22C7# => romdata <= X"C2222010";
    when 16#22C8# => romdata <= X"81C7E008";
    when 16#22C9# => romdata <= X"91E80008";
    when 16#22CA# => romdata <= X"9DE3BFA0";
    when 16#22CB# => romdata <= X"E0066010";
    when 16#22CC# => romdata <= X"2B00003F";
    when 16#22CD# => romdata <= X"A2066014";
    when 16#22CE# => romdata <= X"AA1563FF";
    when 16#22CF# => romdata <= X"A4102000";
    when 16#22D0# => romdata <= X"E8044000";
    when 16#22D1# => romdata <= X"920D0015";
    when 16#22D2# => romdata <= X"400003BC";
    when 16#22D3# => romdata <= X"9010001A";
    when 16#22D4# => romdata <= X"93352010";
    when 16#22D5# => romdata <= X"A606C008";
    when 16#22D6# => romdata <= X"400003B8";
    when 16#22D7# => romdata <= X"9010001A";
    when 16#22D8# => romdata <= X"B734E010";
    when 16#22D9# => romdata <= X"A60CC015";
    when 16#22DA# => romdata <= X"B606C008";
    when 16#22DB# => romdata <= X"832EE010";
    when 16#22DC# => romdata <= X"A6004013";
    when 16#22DD# => romdata <= X"E6244000";
    when 16#22DE# => romdata <= X"A404A001";
    when 16#22DF# => romdata <= X"A2046004";
    when 16#22E0# => romdata <= X"80A40012";
    when 16#22E1# => romdata <= X"14BFFFEF";
    when 16#22E2# => romdata <= X"B736E010";
    when 16#22E3# => romdata <= X"80A6E000";
    when 16#22E4# => romdata <= X"0280000C";
    when 16#22E5# => romdata <= X"01000000";
    when 16#22E6# => romdata <= X"C2066008";
    when 16#22E7# => romdata <= X"80A40001";
    when 16#22E8# => romdata <= X"3680000A";
    when 16#22E9# => romdata <= X"D2066004";
    when 16#22EA# => romdata <= X"82042004";
    when 16#22EB# => romdata <= X"83286002";
    when 16#22EC# => romdata <= X"82064001";
    when 16#22ED# => romdata <= X"A0042001";
    when 16#22EE# => romdata <= X"E0266010";
    when 16#22EF# => romdata <= X"F6206004";
    when 16#22F0# => romdata <= X"81C7E008";
    when 16#22F1# => romdata <= X"91E80019";
    when 16#22F2# => romdata <= X"92026001";
    when 16#22F3# => romdata <= X"7FFFFE16";
    when 16#22F4# => romdata <= X"90100018";
    when 16#22F5# => romdata <= X"D4066010";
    when 16#22F6# => romdata <= X"B4100008";
    when 16#22F7# => romdata <= X"9206600C";
    when 16#22F8# => romdata <= X"9402A002";
    when 16#22F9# => romdata <= X"9002200C";
    when 16#22FA# => romdata <= X"7FFFFC1D";
    when 16#22FB# => romdata <= X"952AA002";
    when 16#22FC# => romdata <= X"C406204C";
    when 16#22FD# => romdata <= X"C2066004";
    when 16#22FE# => romdata <= X"83286002";
    when 16#22FF# => romdata <= X"C6008001";
    when 16#2300# => romdata <= X"C6264000";
    when 16#2301# => romdata <= X"F2208001";
    when 16#2302# => romdata <= X"10BFFFE8";
    when 16#2303# => romdata <= X"B210001A";
    when 16#2304# => romdata <= X"9DE3BFA0";
    when 16#2305# => romdata <= X"828EA003";
    when 16#2306# => romdata <= X"12800032";
    when 16#2307# => romdata <= X"A0100018";
    when 16#2308# => romdata <= X"B53EA002";
    when 16#2309# => romdata <= X"80A6A000";
    when 16#230A# => romdata <= X"02800025";
    when 16#230B# => romdata <= X"01000000";
    when 16#230C# => romdata <= X"E2042048";
    when 16#230D# => romdata <= X"80A46000";
    when 16#230E# => romdata <= X"02800035";
    when 16#230F# => romdata <= X"90100010";
    when 16#2310# => romdata <= X"808EA001";
    when 16#2311# => romdata <= X"1280000F";
    when 16#2312# => romdata <= X"92100019";
    when 16#2313# => romdata <= X"B53EA001";
    when 16#2314# => romdata <= X"80A6A000";
    when 16#2315# => romdata <= X"0280001A";
    when 16#2316# => romdata <= X"01000000";
    when 16#2317# => romdata <= X"D0044000";
    when 16#2318# => romdata <= X"80A22000";
    when 16#2319# => romdata <= X"02800018";
    when 16#231A# => romdata <= X"92100011";
    when 16#231B# => romdata <= X"A2100008";
    when 16#231C# => romdata <= X"808EA001";
    when 16#231D# => romdata <= X"22BFFFF7";
    when 16#231E# => romdata <= X"B53EA001";
    when 16#231F# => romdata <= X"92100019";
    when 16#2320# => romdata <= X"94100011";
    when 16#2321# => romdata <= X"7FFFFF18";
    when 16#2322# => romdata <= X"90100010";
    when 16#2323# => romdata <= X"80A66000";
    when 16#2324# => romdata <= X"02800008";
    when 16#2325# => romdata <= X"B53EA001";
    when 16#2326# => romdata <= X"C404204C";
    when 16#2327# => romdata <= X"C2066004";
    when 16#2328# => romdata <= X"83286002";
    when 16#2329# => romdata <= X"C6008001";
    when 16#232A# => romdata <= X"C6264000";
    when 16#232B# => romdata <= X"F2208001";
    when 16#232C# => romdata <= X"80A6A000";
    when 16#232D# => romdata <= X"12BFFFEA";
    when 16#232E# => romdata <= X"B2100008";
    when 16#232F# => romdata <= X"81C7E008";
    when 16#2330# => romdata <= X"91E80019";
    when 16#2331# => romdata <= X"94100011";
    when 16#2332# => romdata <= X"7FFFFF07";
    when 16#2333# => romdata <= X"90100010";
    when 16#2334# => romdata <= X"D0244000";
    when 16#2335# => romdata <= X"C0220000";
    when 16#2336# => romdata <= X"10BFFFE6";
    when 16#2337# => romdata <= X"A2100008";
    when 16#2338# => romdata <= X"82007FFF";
    when 16#2339# => romdata <= X"05100032";
    when 16#233A# => romdata <= X"83286002";
    when 16#233B# => romdata <= X"8410A268";
    when 16#233C# => romdata <= X"D4008001";
    when 16#233D# => romdata <= X"92100019";
    when 16#233E# => romdata <= X"90100018";
    when 16#233F# => romdata <= X"7FFFFF8B";
    when 16#2340# => romdata <= X"96102000";
    when 16#2341# => romdata <= X"10BFFFC7";
    when 16#2342# => romdata <= X"B2100008";
    when 16#2343# => romdata <= X"7FFFFF7E";
    when 16#2344# => romdata <= X"92102271";
    when 16#2345# => romdata <= X"D0242048";
    when 16#2346# => romdata <= X"A2100008";
    when 16#2347# => romdata <= X"10BFFFC9";
    when 16#2348# => romdata <= X"C0220000";
    when 16#2349# => romdata <= X"9DE3BFA0";
    when 16#234A# => romdata <= X"92102009";
    when 16#234B# => romdata <= X"4000037F";
    when 16#234C# => romdata <= X"9006E008";
    when 16#234D# => romdata <= X"A0100018";
    when 16#234E# => romdata <= X"80A22001";
    when 16#234F# => romdata <= X"82102001";
    when 16#2350# => romdata <= X"04800006";
    when 16#2351# => romdata <= X"92102000";
    when 16#2352# => romdata <= X"83286001";
    when 16#2353# => romdata <= X"80A20001";
    when 16#2354# => romdata <= X"14BFFFFE";
    when 16#2355# => romdata <= X"92026001";
    when 16#2356# => romdata <= X"7FFFFDB3";
    when 16#2357# => romdata <= X"90100010";
    when 16#2358# => romdata <= X"82102001";
    when 16#2359# => romdata <= X"F8222014";
    when 16#235A# => romdata <= X"C2222010";
    when 16#235B# => romdata <= X"80A6A009";
    when 16#235C# => romdata <= X"A406600A";
    when 16#235D# => romdata <= X"04800010";
    when 16#235E# => romdata <= X"A2102009";
    when 16#235F# => romdata <= X"A4066009";
    when 16#2360# => romdata <= X"D64E4011";
    when 16#2361# => romdata <= X"92100008";
    when 16#2362# => romdata <= X"9602FFD0";
    when 16#2363# => romdata <= X"90100010";
    when 16#2364# => romdata <= X"7FFFFF66";
    when 16#2365# => romdata <= X"9410200A";
    when 16#2366# => romdata <= X"A2046001";
    when 16#2367# => romdata <= X"80A68011";
    when 16#2368# => romdata <= X"34BFFFF9";
    when 16#2369# => romdata <= X"D64E4011";
    when 16#236A# => romdata <= X"A404801A";
    when 16#236B# => romdata <= X"A210001A";
    when 16#236C# => romdata <= X"A404BFF8";
    when 16#236D# => romdata <= X"80A6C011";
    when 16#236E# => romdata <= X"0480000D";
    when 16#236F# => romdata <= X"B4102000";
    when 16#2370# => romdata <= X"D64C801A";
    when 16#2371# => romdata <= X"92100008";
    when 16#2372# => romdata <= X"9602FFD0";
    when 16#2373# => romdata <= X"90100010";
    when 16#2374# => romdata <= X"7FFFFF56";
    when 16#2375# => romdata <= X"9410200A";
    when 16#2376# => romdata <= X"B406A001";
    when 16#2377# => romdata <= X"82068011";
    when 16#2378# => romdata <= X"80A6C001";
    when 16#2379# => romdata <= X"34BFFFF8";
    when 16#237A# => romdata <= X"D64C801A";
    when 16#237B# => romdata <= X"81C7E008";
    when 16#237C# => romdata <= X"91E80008";
    when 16#237D# => romdata <= X"9DE3BFA0";
    when 16#237E# => romdata <= X"80A66000";
    when 16#237F# => romdata <= X"12800004";
    when 16#2380# => romdata <= X"A0100018";
    when 16#2381# => romdata <= X"7FFFE6A8";
    when 16#2382# => romdata <= X"93E8001A";
    when 16#2383# => romdata <= X"7FFFE862";
    when 16#2384# => romdata <= X"90100018";
    when 16#2385# => romdata <= X"AC067FF8";
    when 16#2386# => romdata <= X"C405A004";
    when 16#2387# => romdata <= X"A206A00B";
    when 16#2388# => romdata <= X"80A46016";
    when 16#2389# => romdata <= X"18800009";
    when 16#238A# => romdata <= X"82100002";
    when 16#238B# => romdata <= X"A2102010";
    when 16#238C# => romdata <= X"88102000";
    when 16#238D# => romdata <= X"80A4401A";
    when 16#238E# => romdata <= X"1A800009";
    when 16#238F# => romdata <= X"86102010";
    when 16#2390# => romdata <= X"81C7E008";
    when 16#2391# => romdata <= X"91E82000";
    when 16#2392# => romdata <= X"A20C7FF8";
    when 16#2393# => romdata <= X"86100011";
    when 16#2394# => romdata <= X"80A4401A";
    when 16#2395# => romdata <= X"0ABFFFFB";
    when 16#2396# => romdata <= X"8934601F";
    when 16#2397# => romdata <= X"808920FF";
    when 16#2398# => romdata <= X"12BFFFF8";
    when 16#2399# => romdata <= X"AE08BFFC";
    when 16#239A# => romdata <= X"80A5C003";
    when 16#239B# => romdata <= X"16800054";
    when 16#239C# => romdata <= X"A4100017";
    when 16#239D# => romdata <= X"29100034";
    when 16#239E# => romdata <= X"A8152020";
    when 16#239F# => romdata <= X"C8052008";
    when 16#23A0# => romdata <= X"82058017";
    when 16#23A1# => romdata <= X"80A10001";
    when 16#23A2# => romdata <= X"228000F5";
    when 16#23A3# => romdata <= X"82046010";
    when 16#23A4# => romdata <= X"EA006004";
    when 16#23A5# => romdata <= X"9A0D7FFE";
    when 16#23A6# => romdata <= X"9A00400D";
    when 16#23A7# => romdata <= X"DA036004";
    when 16#23A8# => romdata <= X"808B6001";
    when 16#23A9# => romdata <= X"32800064";
    when 16#23AA# => romdata <= X"AA102000";
    when 16#23AB# => romdata <= X"AA0D7FFC";
    when 16#23AC# => romdata <= X"A4054017";
    when 16#23AD# => romdata <= X"80A48003";
    when 16#23AE# => romdata <= X"36800061";
    when 16#23AF# => romdata <= X"C8006008";
    when 16#23B0# => romdata <= X"8088A001";
    when 16#23B1# => romdata <= X"128000A0";
    when 16#23B2# => romdata <= X"80A06000";
    when 16#23B3# => romdata <= X"E6067FF8";
    when 16#23B4# => romdata <= X"A6258013";
    when 16#23B5# => romdata <= X"E404E004";
    when 16#23B6# => romdata <= X"028000F8";
    when 16#23B7# => romdata <= X"A40CBFFC";
    when 16#23B8# => romdata <= X"80A04004";
    when 16#23B9# => romdata <= X"0280005D";
    when 16#23BA# => romdata <= X"84048017";
    when 16#23BB# => romdata <= X"A4054002";
    when 16#23BC# => romdata <= X"80A48003";
    when 16#23BD# => romdata <= X"368000C9";
    when 16#23BE# => romdata <= X"C4006008";
    when 16#23BF# => romdata <= X"A4100002";
    when 16#23C0# => romdata <= X"80A48003";
    when 16#23C1# => romdata <= X"06800091";
    when 16#23C2# => romdata <= X"9210001A";
    when 16#23C3# => romdata <= X"C404E00C";
    when 16#23C4# => romdata <= X"C204E008";
    when 16#23C5# => romdata <= X"9405FFFC";
    when 16#23C6# => romdata <= X"9004E008";
    when 16#23C7# => romdata <= X"C220A008";
    when 16#23C8# => romdata <= X"80A2A024";
    when 16#23C9# => romdata <= X"188000C8";
    when 16#23CA# => romdata <= X"C420600C";
    when 16#23CB# => romdata <= X"80A2A013";
    when 16#23CC# => romdata <= X"82100019";
    when 16#23CD# => romdata <= X"08800018";
    when 16#23CE# => romdata <= X"86100008";
    when 16#23CF# => romdata <= X"C4064000";
    when 16#23D0# => romdata <= X"C424E008";
    when 16#23D1# => romdata <= X"80A2A01B";
    when 16#23D2# => romdata <= X"8604E010";
    when 16#23D3# => romdata <= X"C4066004";
    when 16#23D4# => romdata <= X"C424E00C";
    when 16#23D5# => romdata <= X"08800010";
    when 16#23D6# => romdata <= X"82066008";
    when 16#23D7# => romdata <= X"C4066008";
    when 16#23D8# => romdata <= X"C424E010";
    when 16#23D9# => romdata <= X"80A2A024";
    when 16#23DA# => romdata <= X"8604E018";
    when 16#23DB# => romdata <= X"C4006004";
    when 16#23DC# => romdata <= X"C424E014";
    when 16#23DD# => romdata <= X"12800008";
    when 16#23DE# => romdata <= X"82006008";
    when 16#23DF# => romdata <= X"C4004000";
    when 16#23E0# => romdata <= X"C424E018";
    when 16#23E1# => romdata <= X"8604E020";
    when 16#23E2# => romdata <= X"C4006004";
    when 16#23E3# => romdata <= X"C424E01C";
    when 16#23E4# => romdata <= X"82006008";
    when 16#23E5# => romdata <= X"C4004000";
    when 16#23E6# => romdata <= X"C420C000";
    when 16#23E7# => romdata <= X"B0100008";
    when 16#23E8# => romdata <= X"84100013";
    when 16#23E9# => romdata <= X"C8006004";
    when 16#23EA# => romdata <= X"C820E004";
    when 16#23EB# => romdata <= X"C2006008";
    when 16#23EC# => romdata <= X"C220E008";
    when 16#23ED# => romdata <= X"10800004";
    when 16#23EE# => romdata <= X"C204E004";
    when 16#23EF# => romdata <= X"84100016";
    when 16#23F0# => romdata <= X"B005A008";
    when 16#23F1# => romdata <= X"86248011";
    when 16#23F2# => romdata <= X"80A0E00F";
    when 16#23F3# => romdata <= X"1880000D";
    when 16#23F4# => romdata <= X"92008011";
    when 16#23F5# => romdata <= X"82086001";
    when 16#23F6# => romdata <= X"82104012";
    when 16#23F7# => romdata <= X"C220A004";
    when 16#23F8# => romdata <= X"A4008012";
    when 16#23F9# => romdata <= X"C204A004";
    when 16#23FA# => romdata <= X"82106001";
    when 16#23FB# => romdata <= X"C224A004";
    when 16#23FC# => romdata <= X"7FFFE7E3";
    when 16#23FD# => romdata <= X"90100010";
    when 16#23FE# => romdata <= X"81C7E008";
    when 16#23FF# => romdata <= X"81E80000";
    when 16#2400# => romdata <= X"82086001";
    when 16#2401# => romdata <= X"A2104011";
    when 16#2402# => romdata <= X"E220A004";
    when 16#2403# => romdata <= X"8210E001";
    when 16#2404# => romdata <= X"C2226004";
    when 16#2405# => romdata <= X"82024003";
    when 16#2406# => romdata <= X"90100010";
    when 16#2407# => romdata <= X"C4006004";
    when 16#2408# => romdata <= X"8410A001";
    when 16#2409# => romdata <= X"C4206004";
    when 16#240A# => romdata <= X"7FFFF82D";
    when 16#240B# => romdata <= X"92026008";
    when 16#240C# => romdata <= X"30BFFFF0";
    when 16#240D# => romdata <= X"10BFFFA3";
    when 16#240E# => romdata <= X"82102000";
    when 16#240F# => romdata <= X"C600600C";
    when 16#2410# => romdata <= X"B005A008";
    when 16#2411# => romdata <= X"82100002";
    when 16#2412# => romdata <= X"C621200C";
    when 16#2413# => romdata <= X"84100016";
    when 16#2414# => romdata <= X"10BFFFDD";
    when 16#2415# => romdata <= X"C820E008";
    when 16#2416# => romdata <= X"A4048017";
    when 16#2417# => romdata <= X"82046010";
    when 16#2418# => romdata <= X"AA054012";
    when 16#2419# => romdata <= X"80A54001";
    when 16#241A# => romdata <= X"06BFFFA7";
    when 16#241B# => romdata <= X"80A48003";
    when 16#241C# => romdata <= X"C404E00C";
    when 16#241D# => romdata <= X"C204E008";
    when 16#241E# => romdata <= X"9405FFFC";
    when 16#241F# => romdata <= X"B004E008";
    when 16#2420# => romdata <= X"C220A008";
    when 16#2421# => romdata <= X"80A2A024";
    when 16#2422# => romdata <= X"18800094";
    when 16#2423# => romdata <= X"C420600C";
    when 16#2424# => romdata <= X"80A2A013";
    when 16#2425# => romdata <= X"82100019";
    when 16#2426# => romdata <= X"08800018";
    when 16#2427# => romdata <= X"84100018";
    when 16#2428# => romdata <= X"C4064000";
    when 16#2429# => romdata <= X"C424E008";
    when 16#242A# => romdata <= X"80A2A01B";
    when 16#242B# => romdata <= X"8404E010";
    when 16#242C# => romdata <= X"C6066004";
    when 16#242D# => romdata <= X"C624E00C";
    when 16#242E# => romdata <= X"08800010";
    when 16#242F# => romdata <= X"82066008";
    when 16#2430# => romdata <= X"C4066008";
    when 16#2431# => romdata <= X"C424E010";
    when 16#2432# => romdata <= X"80A2A024";
    when 16#2433# => romdata <= X"8404E018";
    when 16#2434# => romdata <= X"C6006004";
    when 16#2435# => romdata <= X"C624E014";
    when 16#2436# => romdata <= X"12800008";
    when 16#2437# => romdata <= X"82006008";
    when 16#2438# => romdata <= X"C4004000";
    when 16#2439# => romdata <= X"C424E018";
    when 16#243A# => romdata <= X"8404E020";
    when 16#243B# => romdata <= X"C6006004";
    when 16#243C# => romdata <= X"C624E01C";
    when 16#243D# => romdata <= X"82006008";
    when 16#243E# => romdata <= X"C6004000";
    when 16#243F# => romdata <= X"C6208000";
    when 16#2440# => romdata <= X"C6006004";
    when 16#2441# => romdata <= X"C620A004";
    when 16#2442# => romdata <= X"C2006008";
    when 16#2443# => romdata <= X"C220A008";
    when 16#2444# => romdata <= X"8204C011";
    when 16#2445# => romdata <= X"84254011";
    when 16#2446# => romdata <= X"8410A001";
    when 16#2447# => romdata <= X"C4206004";
    when 16#2448# => romdata <= X"C2252008";
    when 16#2449# => romdata <= X"90100010";
    when 16#244A# => romdata <= X"C204E004";
    when 16#244B# => romdata <= X"82086001";
    when 16#244C# => romdata <= X"A2144001";
    when 16#244D# => romdata <= X"7FFFE792";
    when 16#244E# => romdata <= X"E224E004";
    when 16#244F# => romdata <= X"81C7E008";
    when 16#2450# => romdata <= X"81E80000";
    when 16#2451# => romdata <= X"9210001A";
    when 16#2452# => romdata <= X"7FFFE5D7";
    when 16#2453# => romdata <= X"90100010";
    when 16#2454# => romdata <= X"B0922000";
    when 16#2455# => romdata <= X"0280002D";
    when 16#2456# => romdata <= X"84063FF8";
    when 16#2457# => romdata <= X"C205A004";
    when 16#2458# => romdata <= X"86087FFE";
    when 16#2459# => romdata <= X"86058003";
    when 16#245A# => romdata <= X"80A08003";
    when 16#245B# => romdata <= X"02800055";
    when 16#245C# => romdata <= X"9405FFFC";
    when 16#245D# => romdata <= X"80A2A024";
    when 16#245E# => romdata <= X"1880004C";
    when 16#245F# => romdata <= X"80A2A013";
    when 16#2460# => romdata <= X"84100019";
    when 16#2461# => romdata <= X"08800018";
    when 16#2462# => romdata <= X"82100018";
    when 16#2463# => romdata <= X"C2064000";
    when 16#2464# => romdata <= X"C2260000";
    when 16#2465# => romdata <= X"80A2A01B";
    when 16#2466# => romdata <= X"82062008";
    when 16#2467# => romdata <= X"C4066004";
    when 16#2468# => romdata <= X"C4262004";
    when 16#2469# => romdata <= X"08800010";
    when 16#246A# => romdata <= X"84066008";
    when 16#246B# => romdata <= X"C2066008";
    when 16#246C# => romdata <= X"C2262008";
    when 16#246D# => romdata <= X"80A2A024";
    when 16#246E# => romdata <= X"82062010";
    when 16#246F# => romdata <= X"C406600C";
    when 16#2470# => romdata <= X"C426200C";
    when 16#2471# => romdata <= X"12800008";
    when 16#2472# => romdata <= X"84066010";
    when 16#2473# => romdata <= X"C2066010";
    when 16#2474# => romdata <= X"C2262010";
    when 16#2475# => romdata <= X"84066018";
    when 16#2476# => romdata <= X"82062018";
    when 16#2477# => romdata <= X"C6066014";
    when 16#2478# => romdata <= X"C6262014";
    when 16#2479# => romdata <= X"C6008000";
    when 16#247A# => romdata <= X"C6204000";
    when 16#247B# => romdata <= X"C600A004";
    when 16#247C# => romdata <= X"C6206004";
    when 16#247D# => romdata <= X"C400A008";
    when 16#247E# => romdata <= X"C4206008";
    when 16#247F# => romdata <= X"92100019";
    when 16#2480# => romdata <= X"7FFFF7B7";
    when 16#2481# => romdata <= X"90100010";
    when 16#2482# => romdata <= X"7FFFE75D";
    when 16#2483# => romdata <= X"90100010";
    when 16#2484# => romdata <= X"81C7E008";
    when 16#2485# => romdata <= X"81E80000";
    when 16#2486# => romdata <= X"C200600C";
    when 16#2487# => romdata <= X"9405FFFC";
    when 16#2488# => romdata <= X"9004E008";
    when 16#2489# => romdata <= X"C220A00C";
    when 16#248A# => romdata <= X"C4206008";
    when 16#248B# => romdata <= X"80A2A024";
    when 16#248C# => romdata <= X"C404E00C";
    when 16#248D# => romdata <= X"C204E008";
    when 16#248E# => romdata <= X"C220A008";
    when 16#248F# => romdata <= X"08BFFF3C";
    when 16#2490# => romdata <= X"C420600C";
    when 16#2491# => romdata <= X"92100019";
    when 16#2492# => romdata <= X"7FFFFA85";
    when 16#2493# => romdata <= X"B0100008";
    when 16#2494# => romdata <= X"84100013";
    when 16#2495# => romdata <= X"10BFFF5C";
    when 16#2496# => romdata <= X"C204E004";
    when 16#2497# => romdata <= X"EA012004";
    when 16#2498# => romdata <= X"AA0D7FFC";
    when 16#2499# => romdata <= X"9A054017";
    when 16#249A# => romdata <= X"80A34001";
    when 16#249B# => romdata <= X"06BFFF15";
    when 16#249C# => romdata <= X"82100004";
    when 16#249D# => romdata <= X"82058011";
    when 16#249E# => romdata <= X"84234011";
    when 16#249F# => romdata <= X"8410A001";
    when 16#24A0# => romdata <= X"C4206004";
    when 16#24A1# => romdata <= X"C2252008";
    when 16#24A2# => romdata <= X"90100010";
    when 16#24A3# => romdata <= X"C205A004";
    when 16#24A4# => romdata <= X"82086001";
    when 16#24A5# => romdata <= X"A2144001";
    when 16#24A6# => romdata <= X"7FFFE739";
    when 16#24A7# => romdata <= X"E225A004";
    when 16#24A8# => romdata <= X"81C7E008";
    when 16#24A9# => romdata <= X"91E80019";
    when 16#24AA# => romdata <= X"7FFFFA6D";
    when 16#24AB# => romdata <= X"92100019";
    when 16#24AC# => romdata <= X"10BFFFD4";
    when 16#24AD# => romdata <= X"92100019";
    when 16#24AE# => romdata <= X"10BFFF12";
    when 16#24AF# => romdata <= X"A4048017";
    when 16#24B0# => romdata <= X"E400A004";
    when 16#24B1# => romdata <= X"A40CBFFC";
    when 16#24B2# => romdata <= X"84100016";
    when 16#24B3# => romdata <= X"A4048017";
    when 16#24B4# => romdata <= X"10BFFF3D";
    when 16#24B5# => romdata <= X"B005A008";
    when 16#24B6# => romdata <= X"92100019";
    when 16#24B7# => romdata <= X"7FFFFA60";
    when 16#24B8# => romdata <= X"90100018";
    when 16#24B9# => romdata <= X"10BFFF8C";
    when 16#24BA# => romdata <= X"8204C011";
    when 16#24BB# => romdata <= X"9DE3BFA0";
    when 16#24BC# => romdata <= X"80A62000";
    when 16#24BD# => romdata <= X"0280001F";
    when 16#24BE# => romdata <= X"03100032";
    when 16#24BF# => romdata <= X"E4062148";
    when 16#24C0# => romdata <= X"80A4A000";
    when 16#24C1# => romdata <= X"22800014";
    when 16#24C2# => romdata <= X"C206203C";
    when 16#24C3# => romdata <= X"C204A004";
    when 16#24C4# => romdata <= X"A0807FFF";
    when 16#24C5# => romdata <= X"2C80000C";
    when 16#24C6# => romdata <= X"E4048000";
    when 16#24C7# => romdata <= X"A2006001";
    when 16#24C8# => romdata <= X"A32C6002";
    when 16#24C9# => romdata <= X"A2048011";
    when 16#24CA# => romdata <= X"C2044000";
    when 16#24CB# => romdata <= X"9FC04000";
    when 16#24CC# => romdata <= X"A2047FFC";
    when 16#24CD# => romdata <= X"A0843FFF";
    when 16#24CE# => romdata <= X"3CBFFFFD";
    when 16#24CF# => romdata <= X"C2044000";
    when 16#24D0# => romdata <= X"E4048000";
    when 16#24D1# => romdata <= X"80A4A000";
    when 16#24D2# => romdata <= X"32BFFFF2";
    when 16#24D3# => romdata <= X"C204A004";
    when 16#24D4# => romdata <= X"C206203C";
    when 16#24D5# => romdata <= X"80A06000";
    when 16#24D6# => romdata <= X"02800004";
    when 16#24D7# => romdata <= X"01000000";
    when 16#24D8# => romdata <= X"9FC04000";
    when 16#24D9# => romdata <= X"90100018";
    when 16#24DA# => romdata <= X"81C7E008";
    when 16#24DB# => romdata <= X"81E80000";
    when 16#24DC# => romdata <= X"10BFFFE3";
    when 16#24DD# => romdata <= X"F00062C8";
    when 16#24DE# => romdata <= X"9DE3BFA0";
    when 16#24DF# => romdata <= X"D2064000";
    when 16#24E0# => romdata <= X"80A26000";
    when 16#24E1# => romdata <= X"02800004";
    when 16#24E2# => romdata <= X"01000000";
    when 16#24E3# => romdata <= X"7FFFFFFB";
    when 16#24E4# => romdata <= X"90100018";
    when 16#24E5# => romdata <= X"7FFFF752";
    when 16#24E6# => romdata <= X"81E80000";
    when 16#24E7# => romdata <= X"01000000";
    when 16#24E8# => romdata <= X"9DE3BFA0";
    when 16#24E9# => romdata <= X"03100032";
    when 16#24EA# => romdata <= X"C20062C8";
    when 16#24EB# => romdata <= X"80A60001";
    when 16#24EC# => romdata <= X"02800032";
    when 16#24ED# => romdata <= X"01000000";
    when 16#24EE# => romdata <= X"D206204C";
    when 16#24EF# => romdata <= X"80A26000";
    when 16#24F0# => romdata <= X"22800016";
    when 16#24F1# => romdata <= X"E0062148";
    when 16#24F2# => romdata <= X"A2102000";
    when 16#24F3# => romdata <= X"E0024011";
    when 16#24F4# => romdata <= X"80A42000";
    when 16#24F5# => romdata <= X"2280000B";
    when 16#24F6# => romdata <= X"A2046004";
    when 16#24F7# => romdata <= X"92100010";
    when 16#24F8# => romdata <= X"90100018";
    when 16#24F9# => romdata <= X"7FFFF73E";
    when 16#24FA# => romdata <= X"E0040000";
    when 16#24FB# => romdata <= X"80A42000";
    when 16#24FC# => romdata <= X"12BFFFFC";
    when 16#24FD# => romdata <= X"92100010";
    when 16#24FE# => romdata <= X"D206204C";
    when 16#24FF# => romdata <= X"A2046004";
    when 16#2500# => romdata <= X"80A4603C";
    when 16#2501# => romdata <= X"32BFFFF3";
    when 16#2502# => romdata <= X"E0024011";
    when 16#2503# => romdata <= X"7FFFF734";
    when 16#2504# => romdata <= X"90100018";
    when 16#2505# => romdata <= X"E0062148";
    when 16#2506# => romdata <= X"80A42000";
    when 16#2507# => romdata <= X"2280000E";
    when 16#2508# => romdata <= X"D2062054";
    when 16#2509# => romdata <= X"A206214C";
    when 16#250A# => romdata <= X"80A40011";
    when 16#250B# => romdata <= X"2280000A";
    when 16#250C# => romdata <= X"D2062054";
    when 16#250D# => romdata <= X"92100010";
    when 16#250E# => romdata <= X"90100018";
    when 16#250F# => romdata <= X"7FFFF728";
    when 16#2510# => romdata <= X"E0040000";
    when 16#2511# => romdata <= X"80A44010";
    when 16#2512# => romdata <= X"12BFFFFC";
    when 16#2513# => romdata <= X"92100010";
    when 16#2514# => romdata <= X"D2062054";
    when 16#2515# => romdata <= X"80A26000";
    when 16#2516# => romdata <= X"22800005";
    when 16#2517# => romdata <= X"C2062038";
    when 16#2518# => romdata <= X"7FFFF71F";
    when 16#2519# => romdata <= X"90100018";
    when 16#251A# => romdata <= X"C2062038";
    when 16#251B# => romdata <= X"80A06000";
    when 16#251C# => romdata <= X"32800004";
    when 16#251D# => romdata <= X"C206203C";
    when 16#251E# => romdata <= X"81C7E008";
    when 16#251F# => romdata <= X"81E80000";
    when 16#2520# => romdata <= X"9FC04000";
    when 16#2521# => romdata <= X"90100018";
    when 16#2522# => romdata <= X"F20622E0";
    when 16#2523# => romdata <= X"80A66000";
    when 16#2524# => romdata <= X"02BFFFFA";
    when 16#2525# => romdata <= X"01000000";
    when 16#2526# => romdata <= X"7FFFFFB8";
    when 16#2527# => romdata <= X"81E80000";
    when 16#2528# => romdata <= X"01000000";
    when 16#2529# => romdata <= X"82200009";
    when 16#252A# => romdata <= X"051FFC00";
    when 16#252B# => romdata <= X"82104009";
    when 16#252C# => romdata <= X"09200000";
    when 16#252D# => romdata <= X"8330601F";
    when 16#252E# => romdata <= X"882A0004";
    when 16#252F# => romdata <= X"82104004";
    when 16#2530# => romdata <= X"82208001";
    when 16#2531# => romdata <= X"90200001";
    when 16#2532# => romdata <= X"82120001";
    when 16#2533# => romdata <= X"9138601F";
    when 16#2534# => romdata <= X"81C3E008";
    when 16#2535# => romdata <= X"90022001";
    when 16#2536# => romdata <= X"03200000";
    when 16#2537# => romdata <= X"822A0001";
    when 16#2538# => romdata <= X"90200009";
    when 16#2539# => romdata <= X"90120009";
    when 16#253A# => romdata <= X"9132201F";
    when 16#253B# => romdata <= X"90120001";
    when 16#253C# => romdata <= X"031FFC00";
    when 16#253D# => romdata <= X"90204008";
    when 16#253E# => romdata <= X"81C3E008";
    when 16#253F# => romdata <= X"9132201F";
    when 16#2540# => romdata <= X"D252200E";
    when 16#2541# => romdata <= X"03100032";
    when 16#2542# => romdata <= X"D00062C8";
    when 16#2543# => romdata <= X"8213C000";
    when 16#2544# => romdata <= X"400000A2";
    when 16#2545# => romdata <= X"9E104000";
    when 16#2546# => romdata <= X"01000000";
    when 16#2547# => romdata <= X"9DE3BFA0";
    when 16#2548# => romdata <= X"03100032";
    when 16#2549# => romdata <= X"D256200E";
    when 16#254A# => romdata <= X"D00062C8";
    when 16#254B# => romdata <= X"94100019";
    when 16#254C# => romdata <= X"4000011E";
    when 16#254D# => romdata <= X"9610001A";
    when 16#254E# => romdata <= X"80A23FFF";
    when 16#254F# => romdata <= X"02800008";
    when 16#2550# => romdata <= X"03000004";
    when 16#2551# => romdata <= X"C416200C";
    when 16#2552# => romdata <= X"82108001";
    when 16#2553# => romdata <= X"D0262050";
    when 16#2554# => romdata <= X"C236200C";
    when 16#2555# => romdata <= X"81C7E008";
    when 16#2556# => romdata <= X"91E80008";
    when 16#2557# => romdata <= X"C216200C";
    when 16#2558# => romdata <= X"05000004";
    when 16#2559# => romdata <= X"82284002";
    when 16#255A# => romdata <= X"C236200C";
    when 16#255B# => romdata <= X"81C7E008";
    when 16#255C# => romdata <= X"91E80008";
    when 16#255D# => romdata <= X"9DE3BFA0";
    when 16#255E# => romdata <= X"C216200C";
    when 16#255F# => romdata <= X"A0100018";
    when 16#2560# => romdata <= X"80886100";
    when 16#2561# => romdata <= X"A2100019";
    when 16#2562# => romdata <= X"B610001A";
    when 16#2563# => romdata <= X"02800008";
    when 16#2564# => romdata <= X"25100032";
    when 16#2565# => romdata <= X"D004A2C8";
    when 16#2566# => romdata <= X"D256200E";
    when 16#2567# => romdata <= X"94102000";
    when 16#2568# => romdata <= X"40000102";
    when 16#2569# => romdata <= X"96102002";
    when 16#256A# => romdata <= X"C216200C";
    when 16#256B# => romdata <= X"05000004";
    when 16#256C# => romdata <= X"82284002";
    when 16#256D# => romdata <= X"F004A2C8";
    when 16#256E# => romdata <= X"F254200E";
    when 16#256F# => romdata <= X"C234200C";
    when 16#2570# => romdata <= X"4000003C";
    when 16#2571# => romdata <= X"95E80011";
    when 16#2572# => romdata <= X"01000000";
    when 16#2573# => romdata <= X"9DE3BFA0";
    when 16#2574# => romdata <= X"03100032";
    when 16#2575# => romdata <= X"D256200E";
    when 16#2576# => romdata <= X"D00062C8";
    when 16#2577# => romdata <= X"94100019";
    when 16#2578# => romdata <= X"40000104";
    when 16#2579# => romdata <= X"9610001A";
    when 16#257A# => romdata <= X"80A22000";
    when 16#257B# => romdata <= X"26800007";
    when 16#257C# => romdata <= X"C216200C";
    when 16#257D# => romdata <= X"C2062050";
    when 16#257E# => romdata <= X"82004008";
    when 16#257F# => romdata <= X"C2262050";
    when 16#2580# => romdata <= X"81C7E008";
    when 16#2581# => romdata <= X"91E80008";
    when 16#2582# => romdata <= X"05000004";
    when 16#2583# => romdata <= X"82284002";
    when 16#2584# => romdata <= X"C236200C";
    when 16#2585# => romdata <= X"81C7E008";
    when 16#2586# => romdata <= X"91E80008";
    when 16#2587# => romdata <= X"9DE3BFA0";
    when 16#2588# => romdata <= X"808E2003";
    when 16#2589# => romdata <= X"1280001C";
    when 16#258A# => romdata <= X"82100018";
    when 16#258B# => romdata <= X"C2060000";
    when 16#258C# => romdata <= X"1B3FBFBF";
    when 16#258D# => romdata <= X"9A1362FF";
    when 16#258E# => romdata <= X"8400400D";
    when 16#258F# => romdata <= X"82288001";
    when 16#2590# => romdata <= X"09202020";
    when 16#2591# => romdata <= X"88112080";
    when 16#2592# => romdata <= X"80884004";
    when 16#2593# => romdata <= X"12800012";
    when 16#2594# => romdata <= X"82100018";
    when 16#2595# => romdata <= X"82006004";
    when 16#2596# => romdata <= X"C4004000";
    when 16#2597# => romdata <= X"8600800D";
    when 16#2598# => romdata <= X"8428C002";
    when 16#2599# => romdata <= X"80888004";
    when 16#259A# => romdata <= X"3280000C";
    when 16#259B# => romdata <= X"C4484000";
    when 16#259C# => romdata <= X"82006004";
    when 16#259D# => romdata <= X"C4004000";
    when 16#259E# => romdata <= X"8600800D";
    when 16#259F# => romdata <= X"8428C002";
    when 16#25A0# => romdata <= X"80888004";
    when 16#25A1# => romdata <= X"22BFFFF5";
    when 16#25A2# => romdata <= X"82006004";
    when 16#25A3# => romdata <= X"10800003";
    when 16#25A4# => romdata <= X"C4484000";
    when 16#25A5# => romdata <= X"C4484000";
    when 16#25A6# => romdata <= X"80A0A000";
    when 16#25A7# => romdata <= X"32BFFFFE";
    when 16#25A8# => romdata <= X"82006001";
    when 16#25A9# => romdata <= X"B0204018";
    when 16#25AA# => romdata <= X"81C7E008";
    when 16#25AB# => romdata <= X"81E80000";
    when 16#25AC# => romdata <= X"9DE3BFA0";
    when 16#25AD# => romdata <= X"21100038";
    when 16#25AE# => romdata <= X"90100019";
    when 16#25AF# => romdata <= X"9210001A";
    when 16#25B0# => romdata <= X"C0242260";
    when 16#25B1# => romdata <= X"400002A5";
    when 16#25B2# => romdata <= X"9410001B";
    when 16#25B3# => romdata <= X"80A23FFF";
    when 16#25B4# => romdata <= X"02800004";
    when 16#25B5# => romdata <= X"C2042260";
    when 16#25B6# => romdata <= X"81C7E008";
    when 16#25B7# => romdata <= X"91E80008";
    when 16#25B8# => romdata <= X"80A06000";
    when 16#25B9# => romdata <= X"02BFFFFD";
    when 16#25BA# => romdata <= X"01000000";
    when 16#25BB# => romdata <= X"C2260000";
    when 16#25BC# => romdata <= X"81C7E008";
    when 16#25BD# => romdata <= X"91E80008";
    when 16#25BE# => romdata <= X"9DE3BFA0";
    when 16#25BF# => romdata <= X"92100019";
    when 16#25C0# => romdata <= X"400000CE";
    when 16#25C1# => romdata <= X"9010001A";
    when 16#25C2# => romdata <= X"92100008";
    when 16#25C3# => romdata <= X"7FFFE466";
    when 16#25C4# => romdata <= X"90100018";
    when 16#25C5# => romdata <= X"B0922000";
    when 16#25C6# => romdata <= X"0280001E";
    when 16#25C7# => romdata <= X"01000000";
    when 16#25C8# => romdata <= X"D4063FFC";
    when 16#25C9# => romdata <= X"940ABFFC";
    when 16#25CA# => romdata <= X"9402BFFC";
    when 16#25CB# => romdata <= X"80A2A024";
    when 16#25CC# => romdata <= X"18800016";
    when 16#25CD# => romdata <= X"80A2A013";
    when 16#25CE# => romdata <= X"0880000F";
    when 16#25CF# => romdata <= X"82100018";
    when 16#25D0# => romdata <= X"C0260000";
    when 16#25D1# => romdata <= X"C0262004";
    when 16#25D2# => romdata <= X"80A2A01B";
    when 16#25D3# => romdata <= X"0880000A";
    when 16#25D4# => romdata <= X"82062008";
    when 16#25D5# => romdata <= X"C0262008";
    when 16#25D6# => romdata <= X"C026200C";
    when 16#25D7# => romdata <= X"80A2A024";
    when 16#25D8# => romdata <= X"12800005";
    when 16#25D9# => romdata <= X"82062010";
    when 16#25DA# => romdata <= X"C0262010";
    when 16#25DB# => romdata <= X"C0262014";
    when 16#25DC# => romdata <= X"82062018";
    when 16#25DD# => romdata <= X"C0206008";
    when 16#25DE# => romdata <= X"C0204000";
    when 16#25DF# => romdata <= X"C0206004";
    when 16#25E0# => romdata <= X"81C7E008";
    when 16#25E1# => romdata <= X"81E80000";
    when 16#25E2# => romdata <= X"7FFFF9C8";
    when 16#25E3# => romdata <= X"92102000";
    when 16#25E4# => romdata <= X"81C7E008";
    when 16#25E5# => romdata <= X"81E80000";
    when 16#25E6# => romdata <= X"9DE3BFA0";
    when 16#25E7# => romdata <= X"21100038";
    when 16#25E8# => romdata <= X"90100019";
    when 16#25E9# => romdata <= X"40000237";
    when 16#25EA# => romdata <= X"C0242260";
    when 16#25EB# => romdata <= X"80A23FFF";
    when 16#25EC# => romdata <= X"02800004";
    when 16#25ED# => romdata <= X"C2042260";
    when 16#25EE# => romdata <= X"81C7E008";
    when 16#25EF# => romdata <= X"91E80008";
    when 16#25F0# => romdata <= X"80A06000";
    when 16#25F1# => romdata <= X"02BFFFFD";
    when 16#25F2# => romdata <= X"01000000";
    when 16#25F3# => romdata <= X"C2260000";
    when 16#25F4# => romdata <= X"81C7E008";
    when 16#25F5# => romdata <= X"91E80008";
    when 16#25F6# => romdata <= X"9DE3BFA0";
    when 16#25F7# => romdata <= X"80A66000";
    when 16#25F8# => romdata <= X"0280003E";
    when 16#25F9# => romdata <= X"A0102000";
    when 16#25FA# => romdata <= X"7FFFF55B";
    when 16#25FB# => romdata <= X"A4066058";
    when 16#25FC# => romdata <= X"C216600C";
    when 16#25FD# => romdata <= X"80886200";
    when 16#25FE# => romdata <= X"0280003A";
    when 16#25FF# => romdata <= X"01000000";
    when 16#2600# => romdata <= X"23100032";
    when 16#2601# => romdata <= X"D00462C8";
    when 16#2602# => romdata <= X"80A22000";
    when 16#2603# => romdata <= X"22800007";
    when 16#2604# => romdata <= X"C216600C";
    when 16#2605# => romdata <= X"C2022038";
    when 16#2606# => romdata <= X"80A06000";
    when 16#2607# => romdata <= X"0280003B";
    when 16#2608# => romdata <= X"01000000";
    when 16#2609# => romdata <= X"C216600C";
    when 16#260A# => romdata <= X"83286010";
    when 16#260B# => romdata <= X"80A06000";
    when 16#260C# => romdata <= X"02800030";
    when 16#260D# => romdata <= X"83306010";
    when 16#260E# => romdata <= X"80886008";
    when 16#260F# => romdata <= X"1280003F";
    when 16#2610# => romdata <= X"A0102000";
    when 16#2611# => romdata <= X"C206602C";
    when 16#2612# => romdata <= X"80A06000";
    when 16#2613# => romdata <= X"22800008";
    when 16#2614# => romdata <= X"C216600C";
    when 16#2615# => romdata <= X"9FC04000";
    when 16#2616# => romdata <= X"D006601C";
    when 16#2617# => romdata <= X"80A22000";
    when 16#2618# => romdata <= X"26800002";
    when 16#2619# => romdata <= X"A0103FFF";
    when 16#261A# => romdata <= X"C216600C";
    when 16#261B# => romdata <= X"80886080";
    when 16#261C# => romdata <= X"3280002E";
    when 16#261D# => romdata <= X"D2066010";
    when 16#261E# => romdata <= X"D2066030";
    when 16#261F# => romdata <= X"80A26000";
    when 16#2620# => romdata <= X"02800008";
    when 16#2621# => romdata <= X"82066040";
    when 16#2622# => romdata <= X"80A24001";
    when 16#2623# => romdata <= X"22800005";
    when 16#2624# => romdata <= X"C0266030";
    when 16#2625# => romdata <= X"7FFFF612";
    when 16#2626# => romdata <= X"D00462C8";
    when 16#2627# => romdata <= X"C0266030";
    when 16#2628# => romdata <= X"D2066044";
    when 16#2629# => romdata <= X"80A26000";
    when 16#262A# => romdata <= X"22800006";
    when 16#262B# => romdata <= X"C036600C";
    when 16#262C# => romdata <= X"7FFFF60B";
    when 16#262D# => romdata <= X"D00462C8";
    when 16#262E# => romdata <= X"C0266044";
    when 16#262F# => romdata <= X"C036600C";
    when 16#2630# => romdata <= X"4000048A";
    when 16#2631# => romdata <= X"90100012";
    when 16#2632# => romdata <= X"40000467";
    when 16#2633# => romdata <= X"90100012";
    when 16#2634# => romdata <= X"7FFFF509";
    when 16#2635# => romdata <= X"01000000";
    when 16#2636# => romdata <= X"81C7E008";
    when 16#2637# => romdata <= X"91E80010";
    when 16#2638# => romdata <= X"4000046C";
    when 16#2639# => romdata <= X"90100012";
    when 16#263A# => romdata <= X"10BFFFC7";
    when 16#263B# => romdata <= X"23100032";
    when 16#263C# => romdata <= X"4000047E";
    when 16#263D# => romdata <= X"90100012";
    when 16#263E# => romdata <= X"7FFFF4FF";
    when 16#263F# => romdata <= X"A0102000";
    when 16#2640# => romdata <= X"81C7E008";
    when 16#2641# => romdata <= X"91E80010";
    when 16#2642# => romdata <= X"7FFFF544";
    when 16#2643# => romdata <= X"01000000";
    when 16#2644# => romdata <= X"C216600C";
    when 16#2645# => romdata <= X"83286010";
    when 16#2646# => romdata <= X"80A06000";
    when 16#2647# => romdata <= X"12BFFFC7";
    when 16#2648# => romdata <= X"83306010";
    when 16#2649# => romdata <= X"30BFFFF3";
    when 16#264A# => romdata <= X"7FFFF5ED";
    when 16#264B# => romdata <= X"90100018";
    when 16#264C# => romdata <= X"10BFFFD3";
    when 16#264D# => romdata <= X"D2066030";
    when 16#264E# => romdata <= X"7FFFF483";
    when 16#264F# => romdata <= X"90100019";
    when 16#2650# => romdata <= X"10BFFFC1";
    when 16#2651# => romdata <= X"A0100008";
    when 16#2652# => romdata <= X"92100008";
    when 16#2653# => romdata <= X"03100032";
    when 16#2654# => romdata <= X"D00062C8";
    when 16#2655# => romdata <= X"8213C000";
    when 16#2656# => romdata <= X"7FFFFFA0";
    when 16#2657# => romdata <= X"9E104000";
    when 16#2658# => romdata <= X"01000000";
    when 16#2659# => romdata <= X"9DE3BFA0";
    when 16#265A# => romdata <= X"21100038";
    when 16#265B# => romdata <= X"90100019";
    when 16#265C# => romdata <= X"9210001A";
    when 16#265D# => romdata <= X"400001C5";
    when 16#265E# => romdata <= X"C0242260";
    when 16#265F# => romdata <= X"80A23FFF";
    when 16#2660# => romdata <= X"02800004";
    when 16#2661# => romdata <= X"C2042260";
    when 16#2662# => romdata <= X"81C7E008";
    when 16#2663# => romdata <= X"91E80008";
    when 16#2664# => romdata <= X"80A06000";
    when 16#2665# => romdata <= X"02BFFFFD";
    when 16#2666# => romdata <= X"01000000";
    when 16#2667# => romdata <= X"C2260000";
    when 16#2668# => romdata <= X"81C7E008";
    when 16#2669# => romdata <= X"91E80008";
    when 16#266A# => romdata <= X"9DE3BFA0";
    when 16#266B# => romdata <= X"21100038";
    when 16#266C# => romdata <= X"90100019";
    when 16#266D# => romdata <= X"9210001A";
    when 16#266E# => romdata <= X"C0242260";
    when 16#266F# => romdata <= X"400001BA";
    when 16#2670# => romdata <= X"9410001B";
    when 16#2671# => romdata <= X"80A23FFF";
    when 16#2672# => romdata <= X"02800004";
    when 16#2673# => romdata <= X"C2042260";
    when 16#2674# => romdata <= X"81C7E008";
    when 16#2675# => romdata <= X"91E80008";
    when 16#2676# => romdata <= X"80A06000";
    when 16#2677# => romdata <= X"02BFFFFD";
    when 16#2678# => romdata <= X"01000000";
    when 16#2679# => romdata <= X"C2260000";
    when 16#267A# => romdata <= X"81C7E008";
    when 16#267B# => romdata <= X"91E80008";
    when 16#267C# => romdata <= X"9DE3BFA0";
    when 16#267D# => romdata <= X"21100038";
    when 16#267E# => romdata <= X"90100019";
    when 16#267F# => romdata <= X"9210001A";
    when 16#2680# => romdata <= X"C0242260";
    when 16#2681# => romdata <= X"400001AF";
    when 16#2682# => romdata <= X"9410001B";
    when 16#2683# => romdata <= X"80A23FFF";
    when 16#2684# => romdata <= X"02800004";
    when 16#2685# => romdata <= X"C2042260";
    when 16#2686# => romdata <= X"81C7E008";
    when 16#2687# => romdata <= X"91E80008";
    when 16#2688# => romdata <= X"80A06000";
    when 16#2689# => romdata <= X"02BFFFFD";
    when 16#268A# => romdata <= X"01000000";
    when 16#268B# => romdata <= X"C2260000";
    when 16#268C# => romdata <= X"81C7E008";
    when 16#268D# => romdata <= X"91E80008";
    when 16#268E# => romdata <= X"98120009";
    when 16#268F# => romdata <= X"81820000";
    when 16#2690# => romdata <= X"9AAB2FFF";
    when 16#2691# => romdata <= X"02800025";
    when 16#2692# => romdata <= X"98880000";
    when 16#2693# => romdata <= X"99230009";
    when 16#2694# => romdata <= X"99230009";
    when 16#2695# => romdata <= X"99230009";
    when 16#2696# => romdata <= X"99230009";
    when 16#2697# => romdata <= X"99230009";
    when 16#2698# => romdata <= X"99230009";
    when 16#2699# => romdata <= X"99230009";
    when 16#269A# => romdata <= X"99230009";
    when 16#269B# => romdata <= X"99230009";
    when 16#269C# => romdata <= X"99230009";
    when 16#269D# => romdata <= X"99230009";
    when 16#269E# => romdata <= X"99230009";
    when 16#269F# => romdata <= X"99230009";
    when 16#26A0# => romdata <= X"99230009";
    when 16#26A1# => romdata <= X"99230009";
    when 16#26A2# => romdata <= X"99230009";
    when 16#26A3# => romdata <= X"99230009";
    when 16#26A4# => romdata <= X"99230009";
    when 16#26A5# => romdata <= X"99230009";
    when 16#26A6# => romdata <= X"99230009";
    when 16#26A7# => romdata <= X"99230009";
    when 16#26A8# => romdata <= X"99230009";
    when 16#26A9# => romdata <= X"99230009";
    when 16#26AA# => romdata <= X"99230009";
    when 16#26AB# => romdata <= X"99230009";
    when 16#26AC# => romdata <= X"99230009";
    when 16#26AD# => romdata <= X"99230009";
    when 16#26AE# => romdata <= X"99230009";
    when 16#26AF# => romdata <= X"99230009";
    when 16#26B0# => romdata <= X"99230009";
    when 16#26B1# => romdata <= X"99230009";
    when 16#26B2# => romdata <= X"99230009";
    when 16#26B3# => romdata <= X"99230000";
    when 16#26B4# => romdata <= X"81C3E008";
    when 16#26B5# => romdata <= X"91400000";
    when 16#26B6# => romdata <= X"99230009";
    when 16#26B7# => romdata <= X"99230009";
    when 16#26B8# => romdata <= X"99230009";
    when 16#26B9# => romdata <= X"99230009";
    when 16#26BA# => romdata <= X"99230009";
    when 16#26BB# => romdata <= X"99230009";
    when 16#26BC# => romdata <= X"99230009";
    when 16#26BD# => romdata <= X"99230009";
    when 16#26BE# => romdata <= X"99230009";
    when 16#26BF# => romdata <= X"99230009";
    when 16#26C0# => romdata <= X"99230009";
    when 16#26C1# => romdata <= X"99230009";
    when 16#26C2# => romdata <= X"99230000";
    when 16#26C3# => romdata <= X"9B400000";
    when 16#26C4# => romdata <= X"992B200C";
    when 16#26C5# => romdata <= X"9B336014";
    when 16#26C6# => romdata <= X"81C3E008";
    when 16#26C7# => romdata <= X"9013400C";
    when 16#26C8# => romdata <= X"1080000B";
    when 16#26C9# => romdata <= X"86102000";
    when 16#26CA# => romdata <= X"80924008";
    when 16#26CB# => romdata <= X"16800008";
    when 16#26CC# => romdata <= X"861A4008";
    when 16#26CD# => romdata <= X"80924000";
    when 16#26CE# => romdata <= X"16800004";
    when 16#26CF# => romdata <= X"80920000";
    when 16#26D0# => romdata <= X"16800003";
    when 16#26D1# => romdata <= X"92200009";
    when 16#26D2# => romdata <= X"90200008";
    when 16#26D3# => romdata <= X"9A924000";
    when 16#26D4# => romdata <= X"12800005";
    when 16#26D5# => romdata <= X"96100008";
    when 16#26D6# => romdata <= X"91D02002";
    when 16#26D7# => romdata <= X"81C3E008";
    when 16#26D8# => romdata <= X"90100000";
    when 16#26D9# => romdata <= X"80A2C00D";
    when 16#26DA# => romdata <= X"0A800095";
    when 16#26DB# => romdata <= X"94100000";
    when 16#26DC# => romdata <= X"03020000";
    when 16#26DD# => romdata <= X"80A2C001";
    when 16#26DE# => romdata <= X"0A800028";
    when 16#26DF# => romdata <= X"98100000";
    when 16#26E0# => romdata <= X"80A34001";
    when 16#26E1# => romdata <= X"1A80000D";
    when 16#26E2# => romdata <= X"84102001";
    when 16#26E3# => romdata <= X"9B2B6004";
    when 16#26E4# => romdata <= X"10BFFFFC";
    when 16#26E5# => romdata <= X"98032001";
    when 16#26E6# => romdata <= X"9A83400D";
    when 16#26E7# => romdata <= X"1A800007";
    when 16#26E8# => romdata <= X"8400A001";
    when 16#26E9# => romdata <= X"83286004";
    when 16#26EA# => romdata <= X"9B336001";
    when 16#26EB# => romdata <= X"9A034001";
    when 16#26EC# => romdata <= X"10800007";
    when 16#26ED# => romdata <= X"8420A001";
    when 16#26EE# => romdata <= X"80A3400B";
    when 16#26EF# => romdata <= X"0ABFFFF7";
    when 16#26F0# => romdata <= X"01000000";
    when 16#26F1# => romdata <= X"02800002";
    when 16#26F2# => romdata <= X"01000000";
    when 16#26F3# => romdata <= X"84A0A001";
    when 16#26F4# => romdata <= X"06800076";
    when 16#26F5# => romdata <= X"01000000";
    when 16#26F6# => romdata <= X"9622C00D";
    when 16#26F7# => romdata <= X"94102001";
    when 16#26F8# => romdata <= X"1080000A";
    when 16#26F9# => romdata <= X"01000000";
    when 16#26FA# => romdata <= X"952AA001";
    when 16#26FB# => romdata <= X"06800005";
    when 16#26FC# => romdata <= X"9B336001";
    when 16#26FD# => romdata <= X"9622C00D";
    when 16#26FE# => romdata <= X"10800004";
    when 16#26FF# => romdata <= X"9402A001";
    when 16#2700# => romdata <= X"9602C00D";
    when 16#2701# => romdata <= X"9422A001";
    when 16#2702# => romdata <= X"84A0A001";
    when 16#2703# => romdata <= X"16BFFFF7";
    when 16#2704# => romdata <= X"8092C000";
    when 16#2705# => romdata <= X"30800065";
    when 16#2706# => romdata <= X"9B2B6004";
    when 16#2707# => romdata <= X"80A3400B";
    when 16#2708# => romdata <= X"08BFFFFE";
    when 16#2709# => romdata <= X"98832001";
    when 16#270A# => romdata <= X"02800065";
    when 16#270B# => romdata <= X"98232001";
    when 16#270C# => romdata <= X"8092C000";
    when 16#270D# => romdata <= X"952AA004";
    when 16#270E# => romdata <= X"0680002F";
    when 16#270F# => romdata <= X"9B336001";
    when 16#2710# => romdata <= X"96A2C00D";
    when 16#2711# => romdata <= X"06800017";
    when 16#2712# => romdata <= X"9B336001";
    when 16#2713# => romdata <= X"96A2C00D";
    when 16#2714# => romdata <= X"0680000B";
    when 16#2715# => romdata <= X"9B336001";
    when 16#2716# => romdata <= X"96A2C00D";
    when 16#2717# => romdata <= X"06800005";
    when 16#2718# => romdata <= X"9B336001";
    when 16#2719# => romdata <= X"96A2C00D";
    when 16#271A# => romdata <= X"10800050";
    when 16#271B# => romdata <= X"9402A00F";
    when 16#271C# => romdata <= X"9682C00D";
    when 16#271D# => romdata <= X"1080004D";
    when 16#271E# => romdata <= X"9402A00D";
    when 16#271F# => romdata <= X"9682C00D";
    when 16#2720# => romdata <= X"06800005";
    when 16#2721# => romdata <= X"9B336001";
    when 16#2722# => romdata <= X"96A2C00D";
    when 16#2723# => romdata <= X"10800047";
    when 16#2724# => romdata <= X"9402A00B";
    when 16#2725# => romdata <= X"9682C00D";
    when 16#2726# => romdata <= X"10800044";
    when 16#2727# => romdata <= X"9402A009";
    when 16#2728# => romdata <= X"9682C00D";
    when 16#2729# => romdata <= X"0680000B";
    when 16#272A# => romdata <= X"9B336001";
    when 16#272B# => romdata <= X"96A2C00D";
    when 16#272C# => romdata <= X"06800005";
    when 16#272D# => romdata <= X"9B336001";
    when 16#272E# => romdata <= X"96A2C00D";
    when 16#272F# => romdata <= X"1080003B";
    when 16#2730# => romdata <= X"9402A007";
    when 16#2731# => romdata <= X"9682C00D";
    when 16#2732# => romdata <= X"10800038";
    when 16#2733# => romdata <= X"9402A005";
    when 16#2734# => romdata <= X"9682C00D";
    when 16#2735# => romdata <= X"06800005";
    when 16#2736# => romdata <= X"9B336001";
    when 16#2737# => romdata <= X"96A2C00D";
    when 16#2738# => romdata <= X"10800032";
    when 16#2739# => romdata <= X"9402A003";
    when 16#273A# => romdata <= X"9682C00D";
    when 16#273B# => romdata <= X"1080002F";
    when 16#273C# => romdata <= X"9402A001";
    when 16#273D# => romdata <= X"9682C00D";
    when 16#273E# => romdata <= X"06800017";
    when 16#273F# => romdata <= X"9B336001";
    when 16#2740# => romdata <= X"96A2C00D";
    when 16#2741# => romdata <= X"0680000B";
    when 16#2742# => romdata <= X"9B336001";
    when 16#2743# => romdata <= X"96A2C00D";
    when 16#2744# => romdata <= X"06800005";
    when 16#2745# => romdata <= X"9B336001";
    when 16#2746# => romdata <= X"96A2C00D";
    when 16#2747# => romdata <= X"10800023";
    when 16#2748# => romdata <= X"9402BFFF";
    when 16#2749# => romdata <= X"9682C00D";
    when 16#274A# => romdata <= X"10800020";
    when 16#274B# => romdata <= X"9402BFFD";
    when 16#274C# => romdata <= X"9682C00D";
    when 16#274D# => romdata <= X"06800005";
    when 16#274E# => romdata <= X"9B336001";
    when 16#274F# => romdata <= X"96A2C00D";
    when 16#2750# => romdata <= X"1080001A";
    when 16#2751# => romdata <= X"9402BFFB";
    when 16#2752# => romdata <= X"9682C00D";
    when 16#2753# => romdata <= X"10800017";
    when 16#2754# => romdata <= X"9402BFF9";
    when 16#2755# => romdata <= X"9682C00D";
    when 16#2756# => romdata <= X"0680000B";
    when 16#2757# => romdata <= X"9B336001";
    when 16#2758# => romdata <= X"96A2C00D";
    when 16#2759# => romdata <= X"06800005";
    when 16#275A# => romdata <= X"9B336001";
    when 16#275B# => romdata <= X"96A2C00D";
    when 16#275C# => romdata <= X"1080000E";
    when 16#275D# => romdata <= X"9402BFF7";
    when 16#275E# => romdata <= X"9682C00D";
    when 16#275F# => romdata <= X"1080000B";
    when 16#2760# => romdata <= X"9402BFF5";
    when 16#2761# => romdata <= X"9682C00D";
    when 16#2762# => romdata <= X"06800005";
    when 16#2763# => romdata <= X"9B336001";
    when 16#2764# => romdata <= X"96A2C00D";
    when 16#2765# => romdata <= X"10800005";
    when 16#2766# => romdata <= X"9402BFF3";
    when 16#2767# => romdata <= X"9682C00D";
    when 16#2768# => romdata <= X"10800002";
    when 16#2769# => romdata <= X"9402BFF1";
    when 16#276A# => romdata <= X"98A32001";
    when 16#276B# => romdata <= X"16BFFFA2";
    when 16#276C# => romdata <= X"8092C000";
    when 16#276D# => romdata <= X"26800002";
    when 16#276E# => romdata <= X"9422A001";
    when 16#276F# => romdata <= X"8090C000";
    when 16#2770# => romdata <= X"26800002";
    when 16#2771# => romdata <= X"9420000A";
    when 16#2772# => romdata <= X"81C3E008";
    when 16#2773# => romdata <= X"9010000A";
    when 16#2774# => romdata <= X"1080000B";
    when 16#2775# => romdata <= X"86102000";
    when 16#2776# => romdata <= X"80924008";
    when 16#2777# => romdata <= X"16800008";
    when 16#2778# => romdata <= X"86100008";
    when 16#2779# => romdata <= X"80924000";
    when 16#277A# => romdata <= X"16800004";
    when 16#277B# => romdata <= X"80920000";
    when 16#277C# => romdata <= X"16800003";
    when 16#277D# => romdata <= X"92200009";
    when 16#277E# => romdata <= X"90200008";
    when 16#277F# => romdata <= X"9A924000";
    when 16#2780# => romdata <= X"12800005";
    when 16#2781# => romdata <= X"96100008";
    when 16#2782# => romdata <= X"91D02002";
    when 16#2783# => romdata <= X"81C3E008";
    when 16#2784# => romdata <= X"90100000";
    when 16#2785# => romdata <= X"80A2C00D";
    when 16#2786# => romdata <= X"0A800095";
    when 16#2787# => romdata <= X"94100000";
    when 16#2788# => romdata <= X"03020000";
    when 16#2789# => romdata <= X"80A2C001";
    when 16#278A# => romdata <= X"0A800028";
    when 16#278B# => romdata <= X"98100000";
    when 16#278C# => romdata <= X"80A34001";
    when 16#278D# => romdata <= X"1A80000D";
    when 16#278E# => romdata <= X"84102001";
    when 16#278F# => romdata <= X"9B2B6004";
    when 16#2790# => romdata <= X"10BFFFFC";
    when 16#2791# => romdata <= X"98032001";
    when 16#2792# => romdata <= X"9A83400D";
    when 16#2793# => romdata <= X"1A800007";
    when 16#2794# => romdata <= X"8400A001";
    when 16#2795# => romdata <= X"83286004";
    when 16#2796# => romdata <= X"9B336001";
    when 16#2797# => romdata <= X"9A034001";
    when 16#2798# => romdata <= X"10800007";
    when 16#2799# => romdata <= X"8420A001";
    when 16#279A# => romdata <= X"80A3400B";
    when 16#279B# => romdata <= X"0ABFFFF7";
    when 16#279C# => romdata <= X"01000000";
    when 16#279D# => romdata <= X"02800002";
    when 16#279E# => romdata <= X"01000000";
    when 16#279F# => romdata <= X"84A0A001";
    when 16#27A0# => romdata <= X"06800076";
    when 16#27A1# => romdata <= X"01000000";
    when 16#27A2# => romdata <= X"9622C00D";
    when 16#27A3# => romdata <= X"94102001";
    when 16#27A4# => romdata <= X"1080000A";
    when 16#27A5# => romdata <= X"01000000";
    when 16#27A6# => romdata <= X"952AA001";
    when 16#27A7# => romdata <= X"06800005";
    when 16#27A8# => romdata <= X"9B336001";
    when 16#27A9# => romdata <= X"9622C00D";
    when 16#27AA# => romdata <= X"10800004";
    when 16#27AB# => romdata <= X"9402A001";
    when 16#27AC# => romdata <= X"9602C00D";
    when 16#27AD# => romdata <= X"9422A001";
    when 16#27AE# => romdata <= X"84A0A001";
    when 16#27AF# => romdata <= X"16BFFFF7";
    when 16#27B0# => romdata <= X"8092C000";
    when 16#27B1# => romdata <= X"30800065";
    when 16#27B2# => romdata <= X"9B2B6004";
    when 16#27B3# => romdata <= X"80A3400B";
    when 16#27B4# => romdata <= X"08BFFFFE";
    when 16#27B5# => romdata <= X"98832001";
    when 16#27B6# => romdata <= X"02800065";
    when 16#27B7# => romdata <= X"98232001";
    when 16#27B8# => romdata <= X"8092C000";
    when 16#27B9# => romdata <= X"952AA004";
    when 16#27BA# => romdata <= X"0680002F";
    when 16#27BB# => romdata <= X"9B336001";
    when 16#27BC# => romdata <= X"96A2C00D";
    when 16#27BD# => romdata <= X"06800017";
    when 16#27BE# => romdata <= X"9B336001";
    when 16#27BF# => romdata <= X"96A2C00D";
    when 16#27C0# => romdata <= X"0680000B";
    when 16#27C1# => romdata <= X"9B336001";
    when 16#27C2# => romdata <= X"96A2C00D";
    when 16#27C3# => romdata <= X"06800005";
    when 16#27C4# => romdata <= X"9B336001";
    when 16#27C5# => romdata <= X"96A2C00D";
    when 16#27C6# => romdata <= X"10800050";
    when 16#27C7# => romdata <= X"9402A00F";
    when 16#27C8# => romdata <= X"9682C00D";
    when 16#27C9# => romdata <= X"1080004D";
    when 16#27CA# => romdata <= X"9402A00D";
    when 16#27CB# => romdata <= X"9682C00D";
    when 16#27CC# => romdata <= X"06800005";
    when 16#27CD# => romdata <= X"9B336001";
    when 16#27CE# => romdata <= X"96A2C00D";
    when 16#27CF# => romdata <= X"10800047";
    when 16#27D0# => romdata <= X"9402A00B";
    when 16#27D1# => romdata <= X"9682C00D";
    when 16#27D2# => romdata <= X"10800044";
    when 16#27D3# => romdata <= X"9402A009";
    when 16#27D4# => romdata <= X"9682C00D";
    when 16#27D5# => romdata <= X"0680000B";
    when 16#27D6# => romdata <= X"9B336001";
    when 16#27D7# => romdata <= X"96A2C00D";
    when 16#27D8# => romdata <= X"06800005";
    when 16#27D9# => romdata <= X"9B336001";
    when 16#27DA# => romdata <= X"96A2C00D";
    when 16#27DB# => romdata <= X"1080003B";
    when 16#27DC# => romdata <= X"9402A007";
    when 16#27DD# => romdata <= X"9682C00D";
    when 16#27DE# => romdata <= X"10800038";
    when 16#27DF# => romdata <= X"9402A005";
    when 16#27E0# => romdata <= X"9682C00D";
    when 16#27E1# => romdata <= X"06800005";
    when 16#27E2# => romdata <= X"9B336001";
    when 16#27E3# => romdata <= X"96A2C00D";
    when 16#27E4# => romdata <= X"10800032";
    when 16#27E5# => romdata <= X"9402A003";
    when 16#27E6# => romdata <= X"9682C00D";
    when 16#27E7# => romdata <= X"1080002F";
    when 16#27E8# => romdata <= X"9402A001";
    when 16#27E9# => romdata <= X"9682C00D";
    when 16#27EA# => romdata <= X"06800017";
    when 16#27EB# => romdata <= X"9B336001";
    when 16#27EC# => romdata <= X"96A2C00D";
    when 16#27ED# => romdata <= X"0680000B";
    when 16#27EE# => romdata <= X"9B336001";
    when 16#27EF# => romdata <= X"96A2C00D";
    when 16#27F0# => romdata <= X"06800005";
    when 16#27F1# => romdata <= X"9B336001";
    when 16#27F2# => romdata <= X"96A2C00D";
    when 16#27F3# => romdata <= X"10800023";
    when 16#27F4# => romdata <= X"9402BFFF";
    when 16#27F5# => romdata <= X"9682C00D";
    when 16#27F6# => romdata <= X"10800020";
    when 16#27F7# => romdata <= X"9402BFFD";
    when 16#27F8# => romdata <= X"9682C00D";
    when 16#27F9# => romdata <= X"06800005";
    when 16#27FA# => romdata <= X"9B336001";
    when 16#27FB# => romdata <= X"96A2C00D";
    when 16#27FC# => romdata <= X"1080001A";
    when 16#27FD# => romdata <= X"9402BFFB";
    when 16#27FE# => romdata <= X"9682C00D";
    when 16#27FF# => romdata <= X"10800017";
    when 16#2800# => romdata <= X"9402BFF9";
    when 16#2801# => romdata <= X"9682C00D";
    when 16#2802# => romdata <= X"0680000B";
    when 16#2803# => romdata <= X"9B336001";
    when 16#2804# => romdata <= X"96A2C00D";
    when 16#2805# => romdata <= X"06800005";
    when 16#2806# => romdata <= X"9B336001";
    when 16#2807# => romdata <= X"96A2C00D";
    when 16#2808# => romdata <= X"1080000E";
    when 16#2809# => romdata <= X"9402BFF7";
    when 16#280A# => romdata <= X"9682C00D";
    when 16#280B# => romdata <= X"1080000B";
    when 16#280C# => romdata <= X"9402BFF5";
    when 16#280D# => romdata <= X"9682C00D";
    when 16#280E# => romdata <= X"06800005";
    when 16#280F# => romdata <= X"9B336001";
    when 16#2810# => romdata <= X"96A2C00D";
    when 16#2811# => romdata <= X"10800005";
    when 16#2812# => romdata <= X"9402BFF3";
    when 16#2813# => romdata <= X"9682C00D";
    when 16#2814# => romdata <= X"10800002";
    when 16#2815# => romdata <= X"9402BFF1";
    when 16#2816# => romdata <= X"98A32001";
    when 16#2817# => romdata <= X"16BFFFA2";
    when 16#2818# => romdata <= X"8092C000";
    when 16#2819# => romdata <= X"26800002";
    when 16#281A# => romdata <= X"9602C009";
    when 16#281B# => romdata <= X"8090C000";
    when 16#281C# => romdata <= X"26800002";
    when 16#281D# => romdata <= X"9620000B";
    when 16#281E# => romdata <= X"81C3E008";
    when 16#281F# => romdata <= X"9010000B";
    when 16#2820# => romdata <= X"81C3E008";
    when 16#2821# => romdata <= X"90102000";
    when 16#2822# => romdata <= X"03000008";
    when 16#2823# => romdata <= X"90102000";
    when 16#2824# => romdata <= X"C2326008";
    when 16#2825# => romdata <= X"81C3E008";
    when 16#2826# => romdata <= X"C0226030";
    when 16#2827# => romdata <= X"81C3E008";
    when 16#2828# => romdata <= X"90102001";
    when 16#2829# => romdata <= X"9DE3BFA0";
    when 16#282A# => romdata <= X"40000458";
    when 16#282B# => romdata <= X"B0103FFF";
    when 16#282C# => romdata <= X"8210201D";
    when 16#282D# => romdata <= X"C2220000";
    when 16#282E# => romdata <= X"81C7E008";
    when 16#282F# => romdata <= X"81E80000";
    when 16#2830# => romdata <= X"9DE3BFA0";
    when 16#2831# => romdata <= X"80A6A000";
    when 16#2832# => romdata <= X"14800009";
    when 16#2833# => romdata <= X"B0102000";
    when 16#2834# => romdata <= X"30800011";
    when 16#2835# => romdata <= X"0280000E";
    when 16#2836# => romdata <= X"01000000";
    when 16#2837# => romdata <= X"B0062001";
    when 16#2838# => romdata <= X"80A68018";
    when 16#2839# => romdata <= X"0480000C";
    when 16#283A# => romdata <= X"01000000";
    when 16#283B# => romdata <= X"4000004D";
    when 16#283C# => romdata <= X"01000000";
    when 16#283D# => romdata <= X"D02E4018";
    when 16#283E# => romdata <= X"912A2018";
    when 16#283F# => romdata <= X"913A2018";
    when 16#2840# => romdata <= X"80A2200D";
    when 16#2841# => romdata <= X"12BFFFF4";
    when 16#2842# => romdata <= X"80A2200A";
    when 16#2843# => romdata <= X"81C7E008";
    when 16#2844# => romdata <= X"91EE2001";
    when 16#2845# => romdata <= X"81C7E008";
    when 16#2846# => romdata <= X"81E80000";
    when 16#2847# => romdata <= X"05100038";
    when 16#2848# => romdata <= X"C200A264";
    when 16#2849# => romdata <= X"80A06000";
    when 16#284A# => romdata <= X"22800006";
    when 16#284B# => romdata <= X"03100038";
    when 16#284C# => romdata <= X"90004008";
    when 16#284D# => romdata <= X"D020A264";
    when 16#284E# => romdata <= X"81C3E008";
    when 16#284F# => romdata <= X"90100001";
    when 16#2850# => romdata <= X"82106278";
    when 16#2851# => romdata <= X"90004008";
    when 16#2852# => romdata <= X"C220A264";
    when 16#2853# => romdata <= X"D020A264";
    when 16#2854# => romdata <= X"81C3E008";
    when 16#2855# => romdata <= X"90100001";
    when 16#2856# => romdata <= X"9DE3BFA0";
    when 16#2857# => romdata <= X"80A6A000";
    when 16#2858# => romdata <= X"0480001A";
    when 16#2859# => romdata <= X"A0102000";
    when 16#285A# => romdata <= X"10800009";
    when 16#285B# => romdata <= X"D00E4010";
    when 16#285C# => romdata <= X"40000018";
    when 16#285D# => romdata <= X"913A2018";
    when 16#285E# => romdata <= X"A0042001";
    when 16#285F# => romdata <= X"80A68010";
    when 16#2860# => romdata <= X"04800012";
    when 16#2861# => romdata <= X"01000000";
    when 16#2862# => romdata <= X"D00E4010";
    when 16#2863# => romdata <= X"912A2018";
    when 16#2864# => romdata <= X"833A2018";
    when 16#2865# => romdata <= X"80A0600A";
    when 16#2866# => romdata <= X"12BFFFF6";
    when 16#2867# => romdata <= X"01000000";
    when 16#2868# => romdata <= X"4000000C";
    when 16#2869# => romdata <= X"9010200D";
    when 16#286A# => romdata <= X"D00E4010";
    when 16#286B# => romdata <= X"912A2018";
    when 16#286C# => romdata <= X"40000008";
    when 16#286D# => romdata <= X"913A2018";
    when 16#286E# => romdata <= X"A0042001";
    when 16#286F# => romdata <= X"80A68010";
    when 16#2870# => romdata <= X"34BFFFF3";
    when 16#2871# => romdata <= X"D00E4010";
    when 16#2872# => romdata <= X"81C7E008";
    when 16#2873# => romdata <= X"91E8001A";
    when 16#2874# => romdata <= X"03100035";
    when 16#2875# => romdata <= X"C200620C";
    when 16#2876# => romdata <= X"86006004";
    when 16#2877# => romdata <= X"C400C000";
    when 16#2878# => romdata <= X"8088A004";
    when 16#2879# => romdata <= X"02BFFFFE";
    when 16#287A# => romdata <= X"840A20FF";
    when 16#287B# => romdata <= X"C4204000";
    when 16#287C# => romdata <= X"80A2200A";
    when 16#287D# => romdata <= X"02800004";
    when 16#287E# => romdata <= X"01000000";
    when 16#287F# => romdata <= X"81C3E008";
    when 16#2880# => romdata <= X"01000000";
    when 16#2881# => romdata <= X"C400C000";
    when 16#2882# => romdata <= X"8088A004";
    when 16#2883# => romdata <= X"02BFFFFE";
    when 16#2884# => romdata <= X"8410200D";
    when 16#2885# => romdata <= X"C4204000";
    when 16#2886# => romdata <= X"81C3E008";
    when 16#2887# => romdata <= X"01000000";
    when 16#2888# => romdata <= X"03100035";
    when 16#2889# => romdata <= X"C600620C";
    when 16#288A# => romdata <= X"80A0E000";
    when 16#288B# => romdata <= X"8400E004";
    when 16#288C# => romdata <= X"02800007";
    when 16#288D# => romdata <= X"90102000";
    when 16#288E# => romdata <= X"C2008000";
    when 16#288F# => romdata <= X"80886001";
    when 16#2890# => romdata <= X"02BFFFFE";
    when 16#2891# => romdata <= X"01000000";
    when 16#2892# => romdata <= X"D000C000";
    when 16#2893# => romdata <= X"81C3E008";
    when 16#2894# => romdata <= X"01000000";
    when 16#2895# => romdata <= X"A7500000";
    when 16#2896# => romdata <= X"AE100001";
    when 16#2897# => romdata <= X"8334E001";
    when 16#2898# => romdata <= X"29100035";
    when 16#2899# => romdata <= X"E8052214";
    when 16#289A# => romdata <= X"A92CC014";
    when 16#289B# => romdata <= X"82150001";
    when 16#289C# => romdata <= X"81E00000";
    when 16#289D# => romdata <= X"81904000";
    when 16#289E# => romdata <= X"01000000";
    when 16#289F# => romdata <= X"01000000";
    when 16#28A0# => romdata <= X"01000000";
    when 16#28A1# => romdata <= X"E03BA000";
    when 16#28A2# => romdata <= X"E43BA008";
    when 16#28A3# => romdata <= X"E83BA010";
    when 16#28A4# => romdata <= X"EC3BA018";
    when 16#28A5# => romdata <= X"F03BA020";
    when 16#28A6# => romdata <= X"F43BA028";
    when 16#28A7# => romdata <= X"F83BA030";
    when 16#28A8# => romdata <= X"FC3BA038";
    when 16#28A9# => romdata <= X"81E80000";
    when 16#28AA# => romdata <= X"82100017";
    when 16#28AB# => romdata <= X"81C44000";
    when 16#28AC# => romdata <= X"81CC8000";
    when 16#28AD# => romdata <= X"01000000";
    when 16#28AE# => romdata <= X"01000000";
    when 16#28AF# => romdata <= X"01000000";
    when 16#28B0# => romdata <= X"A7500000";
    when 16#28B1# => romdata <= X"A92CE001";
    when 16#28B2# => romdata <= X"2B100035";
    when 16#28B3# => romdata <= X"EA056214";
    when 16#28B4# => romdata <= X"AB34C015";
    when 16#28B5# => romdata <= X"AA154014";
    when 16#28B6# => romdata <= X"81954000";
    when 16#28B7# => romdata <= X"01000000";
    when 16#28B8# => romdata <= X"01000000";
    when 16#28B9# => romdata <= X"01000000";
    when 16#28BA# => romdata <= X"81E80000";
    when 16#28BB# => romdata <= X"81E80000";
    when 16#28BC# => romdata <= X"E01BA000";
    when 16#28BD# => romdata <= X"E41BA008";
    when 16#28BE# => romdata <= X"E81BA010";
    when 16#28BF# => romdata <= X"EC1BA018";
    when 16#28C0# => romdata <= X"F01BA020";
    when 16#28C1# => romdata <= X"F41BA028";
    when 16#28C2# => romdata <= X"F81BA030";
    when 16#28C3# => romdata <= X"FC1BA038";
    when 16#28C4# => romdata <= X"81E00000";
    when 16#28C5# => romdata <= X"81E00000";
    when 16#28C6# => romdata <= X"81C44000";
    when 16#28C7# => romdata <= X"81CC8000";
    when 16#28C8# => romdata <= X"A7500000";
    when 16#28C9# => romdata <= X"2910002B";
    when 16#28CA# => romdata <= X"ADC52198";
    when 16#28CB# => romdata <= X"01000000";
    when 16#28CC# => romdata <= X"27100035";
    when 16#28CD# => romdata <= X"A614E14C";
    when 16#28CE# => romdata <= X"E024C000";
    when 16#28CF# => romdata <= X"818C2020";
    when 16#28D0# => romdata <= X"01000000";
    when 16#28D1# => romdata <= X"01000000";
    when 16#28D2# => romdata <= X"01000000";
    when 16#28D3# => romdata <= X"9DE3BFA0";
    when 16#28D4# => romdata <= X"9DE3BFA0";
    when 16#28D5# => romdata <= X"9DE3BFA0";
    when 16#28D6# => romdata <= X"9DE3BFA0";
    when 16#28D7# => romdata <= X"9DE3BFA0";
    when 16#28D8# => romdata <= X"9DE3BFA0";
    when 16#28D9# => romdata <= X"9DE3BFA0";
    when 16#28DA# => romdata <= X"81E80000";
    when 16#28DB# => romdata <= X"81E80000";
    when 16#28DC# => romdata <= X"81E80000";
    when 16#28DD# => romdata <= X"81E80000";
    when 16#28DE# => romdata <= X"81E80000";
    when 16#28DF# => romdata <= X"81E80000";
    when 16#28E0# => romdata <= X"81E80000";
    when 16#28E1# => romdata <= X"27100035";
    when 16#28E2# => romdata <= X"A614E14C";
    when 16#28E3# => romdata <= X"C024C000";
    when 16#28E4# => romdata <= X"E203A068";
    when 16#28E5# => romdata <= X"A4046004";
    when 16#28E6# => romdata <= X"E223A064";
    when 16#28E7# => romdata <= X"E423A068";
    when 16#28E8# => romdata <= X"108002A9";
    when 16#28E9# => romdata <= X"AC100000";
    when 16#28EA# => romdata <= X"29100035";
    when 16#28EB# => romdata <= X"A8152130";
    when 16#28EC# => romdata <= X"C2252000";
    when 16#28ED# => romdata <= X"C8252004";
    when 16#28EE# => romdata <= X"E0252010";
    when 16#28EF# => romdata <= X"E2252014";
    when 16#28F0# => romdata <= X"E4252018";
    when 16#28F1# => romdata <= X"E825201C";
    when 16#28F2# => romdata <= X"81E80000";
    when 16#28F3# => romdata <= X"83480000";
    when 16#28F4# => romdata <= X"82106F00";
    when 16#28F5# => romdata <= X"81886020";
    when 16#28F6# => romdata <= X"01000000";
    when 16#28F7# => romdata <= X"01000000";
    when 16#28F8# => romdata <= X"01000000";
    when 16#28F9# => romdata <= X"09100035";
    when 16#28FA# => romdata <= X"C8012214";
    when 16#28FB# => romdata <= X"81E00000";
    when 16#28FC# => romdata <= X"88212001";
    when 16#28FD# => romdata <= X"80A920FF";
    when 16#28FE# => romdata <= X"02800003";
    when 16#28FF# => romdata <= X"01000000";
    when 16#2900# => romdata <= X"01000000";
    when 16#2901# => romdata <= X"80A10000";
    when 16#2902# => romdata <= X"12BFFFF9";
    when 16#2903# => romdata <= X"01000000";
    when 16#2904# => romdata <= X"09100035";
    when 16#2905# => romdata <= X"C8012214";
    when 16#2906# => romdata <= X"81E80000";
    when 16#2907# => romdata <= X"80A920FF";
    when 16#2908# => romdata <= X"02800003";
    when 16#2909# => romdata <= X"01000000";
    when 16#290A# => romdata <= X"01000000";
    when 16#290B# => romdata <= X"88212001";
    when 16#290C# => romdata <= X"80A10000";
    when 16#290D# => romdata <= X"12BFFFF9";
    when 16#290E# => romdata <= X"01000000";
    when 16#290F# => romdata <= X"81E00000";
    when 16#2910# => romdata <= X"29100035";
    when 16#2911# => romdata <= X"A8152130";
    when 16#2912# => romdata <= X"C8052004";
    when 16#2913# => romdata <= X"C2052000";
    when 16#2914# => romdata <= X"E0052010";
    when 16#2915# => romdata <= X"E2052014";
    when 16#2916# => romdata <= X"E4052018";
    when 16#2917# => romdata <= X"C025201C";
    when 16#2918# => romdata <= X"818C2000";
    when 16#2919# => romdata <= X"01000000";
    when 16#291A# => romdata <= X"01000000";
    when 16#291B# => romdata <= X"01000000";
    when 16#291C# => romdata <= X"81C48000";
    when 16#291D# => romdata <= X"81CCA004";
    when 16#291E# => romdata <= X"A0142F00";
    when 16#291F# => romdata <= X"818C0000";
    when 16#2920# => romdata <= X"01000000";
    when 16#2921# => romdata <= X"01000000";
    when 16#2922# => romdata <= X"01000000";
    when 16#2923# => romdata <= X"81C48000";
    when 16#2924# => romdata <= X"81CCA004";
    when 16#2925# => romdata <= X"80A66002";
    when 16#2926# => romdata <= X"12800005";
    when 16#2927# => romdata <= X"A8142F00";
    when 16#2928# => romdata <= X"818D0000";
    when 16#2929# => romdata <= X"B0142020";
    when 16#292A# => romdata <= X"3080001F";
    when 16#292B# => romdata <= X"80A66003";
    when 16#292C# => romdata <= X"12800006";
    when 16#292D# => romdata <= X"A80E2F00";
    when 16#292E# => romdata <= X"AA2C2F00";
    when 16#292F# => romdata <= X"A8154014";
    when 16#2930# => romdata <= X"818D0000";
    when 16#2931# => romdata <= X"30800018";
    when 16#2932# => romdata <= X"80A66004";
    when 16#2933# => romdata <= X"12800008";
    when 16#2934# => romdata <= X"A9480000";
    when 16#2935# => romdata <= X"A8152040";
    when 16#2936# => romdata <= X"818D0000";
    when 16#2937# => romdata <= X"01000000";
    when 16#2938# => romdata <= X"01000000";
    when 16#2939# => romdata <= X"01000000";
    when 16#293A# => romdata <= X"3080000F";
    when 16#293B# => romdata <= X"80A66005";
    when 16#293C# => romdata <= X"12800008";
    when 16#293D# => romdata <= X"A9480000";
    when 16#293E# => romdata <= X"A82D2040";
    when 16#293F# => romdata <= X"818D0000";
    when 16#2940# => romdata <= X"01000000";
    when 16#2941# => romdata <= X"01000000";
    when 16#2942# => romdata <= X"01000000";
    when 16#2943# => romdata <= X"30800006";
    when 16#2944# => romdata <= X"80A66006";
    when 16#2945# => romdata <= X"12800003";
    when 16#2946# => romdata <= X"01000000";
    when 16#2947# => romdata <= X"30BFFFA3";
    when 16#2948# => romdata <= X"91D02000";
    when 16#2949# => romdata <= X"81C48000";
    when 16#294A# => romdata <= X"81CCA004";
    when 16#294B# => romdata <= X"92102003";
    when 16#294C# => romdata <= X"81C3E008";
    when 16#294D# => romdata <= X"91D02002";
    when 16#294E# => romdata <= X"92102002";
    when 16#294F# => romdata <= X"81C3E008";
    when 16#2950# => romdata <= X"91D02002";
    when 16#2951# => romdata <= X"92102006";
    when 16#2952# => romdata <= X"81C3E008";
    when 16#2953# => romdata <= X"91D02002";
    when 16#2954# => romdata <= X"27000004";
    when 16#2955# => romdata <= X"A0140013";
    when 16#2956# => romdata <= X"A6142F00";
    when 16#2957# => romdata <= X"818CE000";
    when 16#2958# => romdata <= X"01000000";
    when 16#2959# => romdata <= X"01000000";
    when 16#295A# => romdata <= X"01000000";
    when 16#295B# => romdata <= X"A7480000";
    when 16#295C# => romdata <= X"29000004";
    when 16#295D# => romdata <= X"A68CC014";
    when 16#295E# => romdata <= X"12800003";
    when 16#295F# => romdata <= X"01000000";
    when 16#2960# => romdata <= X"91D02000";
    when 16#2961# => romdata <= X"29100035";
    when 16#2962# => romdata <= X"A81521F4";
    when 16#2963# => romdata <= X"E8050000";
    when 16#2964# => romdata <= X"2B100035";
    when 16#2965# => romdata <= X"AA1561F0";
    when 16#2966# => romdata <= X"EA054000";
    when 16#2967# => romdata <= X"80A50015";
    when 16#2968# => romdata <= X"0280002D";
    when 16#2969# => romdata <= X"01000000";
    when 16#296A# => romdata <= X"80A00015";
    when 16#296B# => romdata <= X"02800013";
    when 16#296C# => romdata <= X"01000000";
    when 16#296D# => romdata <= X"C13D6000";
    when 16#296E# => romdata <= X"C53D6008";
    when 16#296F# => romdata <= X"C93D6010";
    when 16#2970# => romdata <= X"CD3D6018";
    when 16#2971# => romdata <= X"D13D6020";
    when 16#2972# => romdata <= X"D53D6028";
    when 16#2973# => romdata <= X"D93D6030";
    when 16#2974# => romdata <= X"DD3D6038";
    when 16#2975# => romdata <= X"E13D6040";
    when 16#2976# => romdata <= X"E53D6048";
    when 16#2977# => romdata <= X"E93D6050";
    when 16#2978# => romdata <= X"ED3D6058";
    when 16#2979# => romdata <= X"F13D6060";
    when 16#297A# => romdata <= X"F53D6068";
    when 16#297B# => romdata <= X"F93D6070";
    when 16#297C# => romdata <= X"FD3D6078";
    when 16#297D# => romdata <= X"C12D6080";
    when 16#297E# => romdata <= X"2D100035";
    when 16#297F# => romdata <= X"AC15A1F0";
    when 16#2980# => romdata <= X"E8258000";
    when 16#2981# => romdata <= X"80A00014";
    when 16#2982# => romdata <= X"02800013";
    when 16#2983# => romdata <= X"01000000";
    when 16#2984# => romdata <= X"C11D2000";
    when 16#2985# => romdata <= X"C51D2008";
    when 16#2986# => romdata <= X"C91D2010";
    when 16#2987# => romdata <= X"CD1D2018";
    when 16#2988# => romdata <= X"D11D2020";
    when 16#2989# => romdata <= X"D51D2028";
    when 16#298A# => romdata <= X"D91D2030";
    when 16#298B# => romdata <= X"DD1D2038";
    when 16#298C# => romdata <= X"E11D2040";
    when 16#298D# => romdata <= X"E51D2048";
    when 16#298E# => romdata <= X"E91D2050";
    when 16#298F# => romdata <= X"ED1D2058";
    when 16#2990# => romdata <= X"F11D2060";
    when 16#2991# => romdata <= X"F51D2068";
    when 16#2992# => romdata <= X"F91D2070";
    when 16#2993# => romdata <= X"FD1D2078";
    when 16#2994# => romdata <= X"C10D2080";
    when 16#2995# => romdata <= X"818C2000";
    when 16#2996# => romdata <= X"01000000";
    when 16#2997# => romdata <= X"01000000";
    when 16#2998# => romdata <= X"01000000";
    when 16#2999# => romdata <= X"81C44000";
    when 16#299A# => romdata <= X"81CC8000";
    when 16#299B# => romdata <= X"81C3E008";
    when 16#299C# => romdata <= X"01000000";
    when 16#299D# => romdata <= X"81C3E008";
    when 16#299E# => romdata <= X"01000000";
    when 16#299F# => romdata <= X"81C3E008";
    when 16#29A0# => romdata <= X"01000000";
    when 16#29A1# => romdata <= X"AE25A010";
    when 16#29A2# => romdata <= X"A7500000";
    when 16#29A3# => romdata <= X"2D100029";
    when 16#29A4# => romdata <= X"AC15A298";
    when 16#29A5# => romdata <= X"2910002B";
    when 16#29A6# => romdata <= X"81C52360";
    when 16#29A7# => romdata <= X"01000000";
    when 16#29A8# => romdata <= X"11100035";
    when 16#29A9# => romdata <= X"90122200";
    when 16#29AA# => romdata <= X"D2020000";
    when 16#29AB# => romdata <= X"92026001";
    when 16#29AC# => romdata <= X"D2220000";
    when 16#29AD# => romdata <= X"932DE008";
    when 16#29AE# => romdata <= X"902C2F00";
    when 16#29AF# => romdata <= X"92120009";
    when 16#29B0# => romdata <= X"11100035";
    when 16#29B1# => romdata <= X"901221F8";
    when 16#29B2# => romdata <= X"D0020000";
    when 16#29B3# => romdata <= X"80A00008";
    when 16#29B4# => romdata <= X"22800002";
    when 16#29B5# => romdata <= X"92126F00";
    when 16#29B6# => romdata <= X"818A6020";
    when 16#29B7# => romdata <= X"01000000";
    when 16#29B8# => romdata <= X"01000000";
    when 16#29B9# => romdata <= X"01000000";
    when 16#29BA# => romdata <= X"90100017";
    when 16#29BB# => romdata <= X"40000037";
    when 16#29BC# => romdata <= X"9203A0F8";
    when 16#29BD# => romdata <= X"92142F00";
    when 16#29BE# => romdata <= X"818A6020";
    when 16#29BF# => romdata <= X"01000000";
    when 16#29C0# => romdata <= X"01000000";
    when 16#29C1# => romdata <= X"01000000";
    when 16#29C2# => romdata <= X"11100035";
    when 16#29C3# => romdata <= X"90122200";
    when 16#29C4# => romdata <= X"D2020000";
    when 16#29C5# => romdata <= X"92226001";
    when 16#29C6# => romdata <= X"D2220000";
    when 16#29C7# => romdata <= X"10800239";
    when 16#29C8# => romdata <= X"AC100000";
    when 16#29C9# => romdata <= X"9DE3BFA0";
    when 16#29CA# => romdata <= X"1B100037";
    when 16#29CB# => romdata <= X"892E6002";
    when 16#29CC# => romdata <= X"9A136330";
    when 16#29CD# => romdata <= X"80A6601F";
    when 16#29CE# => romdata <= X"82102000";
    when 16#29CF# => romdata <= X"14800017";
    when 16#29D0# => romdata <= X"C6034004";
    when 16#29D1# => romdata <= X"B32E6004";
    when 16#29D2# => romdata <= X"19100037";
    when 16#29D3# => romdata <= X"80A0E000";
    when 16#29D4# => romdata <= X"981323B0";
    when 16#29D5# => romdata <= X"0280000D";
    when 16#29D6# => romdata <= X"8406400C";
    when 16#29D7# => romdata <= X"80A0C002";
    when 16#29D8# => romdata <= X"12800006";
    when 16#29D9# => romdata <= X"82100003";
    when 16#29DA# => romdata <= X"1080000E";
    when 16#29DB# => romdata <= X"C206400C";
    when 16#29DC# => romdata <= X"2280000C";
    when 16#29DD# => romdata <= X"C206400C";
    when 16#29DE# => romdata <= X"C200600C";
    when 16#29DF# => romdata <= X"80A06000";
    when 16#29E0# => romdata <= X"12BFFFFC";
    when 16#29E1# => romdata <= X"80A08001";
    when 16#29E2# => romdata <= X"C4234004";
    when 16#29E3# => romdata <= X"F026400C";
    when 16#29E4# => romdata <= X"C620A00C";
    when 16#29E5# => romdata <= X"82102000";
    when 16#29E6# => romdata <= X"81C7E008";
    when 16#29E7# => romdata <= X"91E80001";
    when 16#29E8# => romdata <= X"F026400C";
    when 16#29E9# => romdata <= X"81C7E008";
    when 16#29EA# => romdata <= X"91E80001";
    when 16#29EB# => romdata <= X"912A2002";
    when 16#29EC# => romdata <= X"03100037";
    when 16#29ED# => romdata <= X"82106330";
    when 16#29EE# => romdata <= X"C4004008";
    when 16#29EF# => romdata <= X"C422600C";
    when 16#29F0# => romdata <= X"81C3E008";
    when 16#29F1# => romdata <= X"D2204008";
    when 16#29F2# => romdata <= X"9DE3BFA0";
    when 16#29F3# => romdata <= X"05100035";
    when 16#29F4# => romdata <= X"8210A204";
    when 16#29F5# => romdata <= X"C2006004";
    when 16#29F6# => romdata <= X"80A04018";
    when 16#29F7# => romdata <= X"22800040";
    when 16#29F8# => romdata <= X"C400A204";
    when 16#29F9# => romdata <= X"80A62000";
    when 16#29FA# => romdata <= X"22800002";
    when 16#29FB# => romdata <= X"B0100001";
    when 16#29FC# => romdata <= X"A32E2002";
    when 16#29FD# => romdata <= X"03100037";
    when 16#29FE# => romdata <= X"82106330";
    when 16#29FF# => romdata <= X"E0004011";
    when 16#2A00# => romdata <= X"80A42000";
    when 16#2A01# => romdata <= X"02800034";
    when 16#2A02# => romdata <= X"29100038";
    when 16#2A03# => romdata <= X"2D100038";
    when 16#2A04# => romdata <= X"2B100038";
    when 16#2A05# => romdata <= X"27100038";
    when 16#2A06# => romdata <= X"A81521B0";
    when 16#2A07# => romdata <= X"AC15A234";
    when 16#2A08# => romdata <= X"AA156238";
    when 16#2A09# => romdata <= X"1080001D";
    when 16#2A0A# => romdata <= X"A614E1B4";
    when 16#2A0B# => romdata <= X"A4100013";
    when 16#2A0C# => romdata <= X"8400A001";
    when 16#2A0D# => romdata <= X"C4248011";
    when 16#2A0E# => romdata <= X"C4058000";
    when 16#2A0F# => romdata <= X"80A0A000";
    when 16#2A10# => romdata <= X"22800006";
    when 16#2A11# => romdata <= X"D2042008";
    when 16#2A12# => romdata <= X"9FC08000";
    when 16#2A13# => romdata <= X"01000000";
    when 16#2A14# => romdata <= X"C2040000";
    when 16#2A15# => romdata <= X"D2042008";
    when 16#2A16# => romdata <= X"90100018";
    when 16#2A17# => romdata <= X"9FC04000";
    when 16#2A18# => romdata <= X"94100019";
    when 16#2A19# => romdata <= X"C2054000";
    when 16#2A1A# => romdata <= X"80A06000";
    when 16#2A1B# => romdata <= X"22800005";
    when 16#2A1C# => romdata <= X"C2048011";
    when 16#2A1D# => romdata <= X"9FC04000";
    when 16#2A1E# => romdata <= X"01000000";
    when 16#2A1F# => romdata <= X"C2048011";
    when 16#2A20# => romdata <= X"82007FFF";
    when 16#2A21# => romdata <= X"C2248011";
    when 16#2A22# => romdata <= X"E004200C";
    when 16#2A23# => romdata <= X"80A42000";
    when 16#2A24# => romdata <= X"02800011";
    when 16#2A25# => romdata <= X"01000000";
    when 16#2A26# => romdata <= X"C2040000";
    when 16#2A27# => romdata <= X"80A06000";
    when 16#2A28# => romdata <= X"22BFFFFB";
    when 16#2A29# => romdata <= X"E004200C";
    when 16#2A2A# => romdata <= X"C4050000";
    when 16#2A2B# => romdata <= X"80A0A000";
    when 16#2A2C# => romdata <= X"12BFFFDF";
    when 16#2A2D# => romdata <= X"C404C011";
    when 16#2A2E# => romdata <= X"80A0A000";
    when 16#2A2F# => romdata <= X"02BFFFDD";
    when 16#2A30# => romdata <= X"A4100013";
    when 16#2A31# => romdata <= X"E004200C";
    when 16#2A32# => romdata <= X"80A42000";
    when 16#2A33# => romdata <= X"32BFFFF4";
    when 16#2A34# => romdata <= X"C2040000";
    when 16#2A35# => romdata <= X"81C7E008";
    when 16#2A36# => romdata <= X"81E80000";
    when 16#2A37# => romdata <= X"F000A0C0";
    when 16#2A38# => romdata <= X"10BFFFC1";
    when 16#2A39# => romdata <= X"B00E201F";
    when 16#2A3A# => romdata <= X"8C10000F";
    when 16#2A3B# => romdata <= X"A7480000";
    when 16#2A3C# => romdata <= X"8B34E018";
    when 16#2A3D# => romdata <= X"8A09600F";
    when 16#2A3E# => romdata <= X"80A16003";
    when 16#2A3F# => romdata <= X"0280000C";
    when 16#2A40# => romdata <= X"0B100035";
    when 16#2A41# => romdata <= X"8A11620C";
    when 16#2A42# => romdata <= X"09200000";
    when 16#2A43# => romdata <= X"88112070";
    when 16#2A44# => romdata <= X"C8214000";
    when 16#2A45# => romdata <= X"0B100035";
    when 16#2A46# => romdata <= X"8A116228";
    when 16#2A47# => romdata <= X"09200000";
    when 16#2A48# => romdata <= X"88112040";
    when 16#2A49# => romdata <= X"C8214000";
    when 16#2A4A# => romdata <= X"10800039";
    when 16#2A4B# => romdata <= X"90102001";
    when 16#2A4C# => romdata <= X"92102006";
    when 16#2A4D# => romdata <= X"400001FC";
    when 16#2A4E# => romdata <= X"01000000";
    when 16#2A4F# => romdata <= X"80A00008";
    when 16#2A50# => romdata <= X"02800033";
    when 16#2A51# => romdata <= X"01000000";
    when 16#2A52# => romdata <= X"C2022010";
    when 16#2A53# => romdata <= X"113FFC00";
    when 16#2A54# => romdata <= X"82084008";
    when 16#2A55# => romdata <= X"110003FC";
    when 16#2A56# => romdata <= X"84104008";
    when 16#2A57# => romdata <= X"90100002";
    when 16#2A58# => romdata <= X"92102001";
    when 16#2A59# => romdata <= X"9410200C";
    when 16#2A5A# => romdata <= X"40000205";
    when 16#2A5B# => romdata <= X"01000000";
    when 16#2A5C# => romdata <= X"80A00008";
    when 16#2A5D# => romdata <= X"02800026";
    when 16#2A5E# => romdata <= X"01000000";
    when 16#2A5F# => romdata <= X"40000215";
    when 16#2A60# => romdata <= X"92100001";
    when 16#2A61# => romdata <= X"0B100035";
    when 16#2A62# => romdata <= X"8A11620C";
    when 16#2A63# => romdata <= X"D2214000";
    when 16#2A64# => romdata <= X"90100002";
    when 16#2A65# => romdata <= X"92102001";
    when 16#2A66# => romdata <= X"94102011";
    when 16#2A67# => romdata <= X"400001F8";
    when 16#2A68# => romdata <= X"01000000";
    when 16#2A69# => romdata <= X"80A00008";
    when 16#2A6A# => romdata <= X"02800019";
    when 16#2A6B# => romdata <= X"01000000";
    when 16#2A6C# => romdata <= X"40000208";
    when 16#2A6D# => romdata <= X"92100001";
    when 16#2A6E# => romdata <= X"92026010";
    when 16#2A6F# => romdata <= X"0B100035";
    when 16#2A70# => romdata <= X"8A116228";
    when 16#2A71# => romdata <= X"D2214000";
    when 16#2A72# => romdata <= X"90100002";
    when 16#2A73# => romdata <= X"92102001";
    when 16#2A74# => romdata <= X"9410200D";
    when 16#2A75# => romdata <= X"400001EA";
    when 16#2A76# => romdata <= X"01000000";
    when 16#2A77# => romdata <= X"80A00008";
    when 16#2A78# => romdata <= X"0280000B";
    when 16#2A79# => romdata <= X"01000000";
    when 16#2A7A# => romdata <= X"400001FA";
    when 16#2A7B# => romdata <= X"92100001";
    when 16#2A7C# => romdata <= X"0B100035";
    when 16#2A7D# => romdata <= X"8A116204";
    when 16#2A7E# => romdata <= X"D2214000";
    when 16#2A7F# => romdata <= X"D4026010";
    when 16#2A80# => romdata <= X"9532A010";
    when 16#2A81# => romdata <= X"940AA00F";
    when 16#2A82# => romdata <= X"D4216004";
    when 16#2A83# => romdata <= X"9E100006";
    when 16#2A84# => romdata <= X"81C3E008";
    when 16#2A85# => romdata <= X"01000000";
    when 16#2A86# => romdata <= X"03100035";
    when 16#2A87# => romdata <= X"82106220";
    when 16#2A88# => romdata <= X"82102001";
    when 16#2A89# => romdata <= X"91D02000";
    when 16#2A8A# => romdata <= X"81C3E008";
    when 16#2A8B# => romdata <= X"01000000";
    when 16#2A8C# => romdata <= X"9DE3BFA0";
    when 16#2A8D# => romdata <= X"03100038";
    when 16#2A8E# => romdata <= X"C2006240";
    when 16#2A8F# => romdata <= X"84100018";
    when 16#2A90# => romdata <= X"80A06000";
    when 16#2A91# => romdata <= X"02800006";
    when 16#2A92# => romdata <= X"B0102000";
    when 16#2A93# => romdata <= X"90100002";
    when 16#2A94# => romdata <= X"9FC04000";
    when 16#2A95# => romdata <= X"92100019";
    when 16#2A96# => romdata <= X"B0100008";
    when 16#2A97# => romdata <= X"81C7E008";
    when 16#2A98# => romdata <= X"81E80000";
    when 16#2A99# => romdata <= X"9DE3BFA0";
    when 16#2A9A# => romdata <= X"03100038";
    when 16#2A9B# => romdata <= X"C2006244";
    when 16#2A9C# => romdata <= X"80A06000";
    when 16#2A9D# => romdata <= X"02800005";
    when 16#2A9E# => romdata <= X"84102000";
    when 16#2A9F# => romdata <= X"9FC04000";
    when 16#2AA0# => romdata <= X"90100018";
    when 16#2AA1# => romdata <= X"84100008";
    when 16#2AA2# => romdata <= X"81C7E008";
    when 16#2AA3# => romdata <= X"91E80002";
    when 16#2AA4# => romdata <= X"9DE3BFA0";
    when 16#2AA5# => romdata <= X"03100038";
    when 16#2AA6# => romdata <= X"C200624C";
    when 16#2AA7# => romdata <= X"80A06000";
    when 16#2AA8# => romdata <= X"02800005";
    when 16#2AA9# => romdata <= X"84102000";
    when 16#2AAA# => romdata <= X"9FC04000";
    when 16#2AAB# => romdata <= X"90100018";
    when 16#2AAC# => romdata <= X"84100008";
    when 16#2AAD# => romdata <= X"81C7E008";
    when 16#2AAE# => romdata <= X"91E80002";
    when 16#2AAF# => romdata <= X"9DE3BFA0";
    when 16#2AB0# => romdata <= X"03100038";
    when 16#2AB1# => romdata <= X"C2006248";
    when 16#2AB2# => romdata <= X"80A06000";
    when 16#2AB3# => romdata <= X"02800005";
    when 16#2AB4# => romdata <= X"84102000";
    when 16#2AB5# => romdata <= X"9FC04000";
    when 16#2AB6# => romdata <= X"90100018";
    when 16#2AB7# => romdata <= X"84100008";
    when 16#2AB8# => romdata <= X"81C7E008";
    when 16#2AB9# => romdata <= X"91E80002";
    when 16#2ABA# => romdata <= X"9DE3BFA0";
    when 16#2ABB# => romdata <= X"03100038";
    when 16#2ABC# => romdata <= X"C2006250";
    when 16#2ABD# => romdata <= X"80A06000";
    when 16#2ABE# => romdata <= X"02800005";
    when 16#2ABF# => romdata <= X"84102000";
    when 16#2AC0# => romdata <= X"9FC04000";
    when 16#2AC1# => romdata <= X"90100018";
    when 16#2AC2# => romdata <= X"84100008";
    when 16#2AC3# => romdata <= X"81C7E008";
    when 16#2AC4# => romdata <= X"91E80002";
    when 16#2AC5# => romdata <= X"9DE3BFA0";
    when 16#2AC6# => romdata <= X"03100038";
    when 16#2AC7# => romdata <= X"C2006254";
    when 16#2AC8# => romdata <= X"80A06000";
    when 16#2AC9# => romdata <= X"02800005";
    when 16#2ACA# => romdata <= X"84102000";
    when 16#2ACB# => romdata <= X"9FC04000";
    when 16#2ACC# => romdata <= X"90100018";
    when 16#2ACD# => romdata <= X"84100008";
    when 16#2ACE# => romdata <= X"81C7E008";
    when 16#2ACF# => romdata <= X"91E80002";
    when 16#2AD0# => romdata <= X"9DE3BFA0";
    when 16#2AD1# => romdata <= X"03100038";
    when 16#2AD2# => romdata <= X"C2006258";
    when 16#2AD3# => romdata <= X"80A06000";
    when 16#2AD4# => romdata <= X"02800005";
    when 16#2AD5# => romdata <= X"84102000";
    when 16#2AD6# => romdata <= X"9FC04000";
    when 16#2AD7# => romdata <= X"90100018";
    when 16#2AD8# => romdata <= X"84100008";
    when 16#2AD9# => romdata <= X"81C7E008";
    when 16#2ADA# => romdata <= X"91E80002";
    when 16#2ADB# => romdata <= X"9DE3BFA0";
    when 16#2ADC# => romdata <= X"03100038";
    when 16#2ADD# => romdata <= X"C200625C";
    when 16#2ADE# => romdata <= X"84100018";
    when 16#2ADF# => romdata <= X"80A06000";
    when 16#2AE0# => romdata <= X"02800006";
    when 16#2AE1# => romdata <= X"B0102000";
    when 16#2AE2# => romdata <= X"90100002";
    when 16#2AE3# => romdata <= X"9FC04000";
    when 16#2AE4# => romdata <= X"92100019";
    when 16#2AE5# => romdata <= X"B0100008";
    when 16#2AE6# => romdata <= X"81C7E008";
    when 16#2AE7# => romdata <= X"81E80000";
    when 16#2AE8# => romdata <= X"01000000";
    when 16#2AE9# => romdata <= X"0310002B";
    when 16#2AEA# => romdata <= X"82106070";
    when 16#2AEB# => romdata <= X"9FC04000";
    when 16#2AEC# => romdata <= X"01000000";
    when 16#2AED# => romdata <= X"03100000";
    when 16#2AEE# => romdata <= X"82106000";
    when 16#2AEF# => romdata <= X"81984000";
    when 16#2AF0# => romdata <= X"0310002B";
    when 16#2AF1# => romdata <= X"821060F4";
    when 16#2AF2# => romdata <= X"9FC04000";
    when 16#2AF3# => romdata <= X"01000000";
    when 16#2AF4# => romdata <= X"0310002B";
    when 16#2AF5# => romdata <= X"82106060";
    when 16#2AF6# => romdata <= X"9FC04000";
    when 16#2AF7# => romdata <= X"01000000";
    when 16#2AF8# => romdata <= X"8B480000";
    when 16#2AF9# => romdata <= X"8B316018";
    when 16#2AFA# => romdata <= X"8A096003";
    when 16#2AFB# => romdata <= X"80A16003";
    when 16#2AFC# => romdata <= X"12800007";
    when 16#2AFD# => romdata <= X"01000000";
    when 16#2AFE# => romdata <= X"8B444000";
    when 16#2AFF# => romdata <= X"8B31601C";
    when 16#2B00# => romdata <= X"80A14000";
    when 16#2B01# => romdata <= X"12800006";
    when 16#2B02# => romdata <= X"01000000";
    when 16#2B03# => romdata <= X"7FFFFF37";
    when 16#2B04# => romdata <= X"01000000";
    when 16#2B05# => romdata <= X"7FFFD961";
    when 16#2B06# => romdata <= X"01000000";
    when 16#2B07# => romdata <= X"9C23A040";
    when 16#2B08# => romdata <= X"7FFFD8F8";
    when 16#2B09# => romdata <= X"01000000";
    when 16#2B0A# => romdata <= X"82102001";
    when 16#2B0B# => romdata <= X"91D02000";
    when 16#2B0C# => romdata <= X"01000000";
    when 16#2B0D# => romdata <= X"29000004";
    when 16#2B0E# => romdata <= X"A68C0014";
    when 16#2B0F# => romdata <= X"32800003";
    when 16#2B10# => romdata <= X"A02C0014";
    when 16#2B11# => romdata <= X"91D02000";
    when 16#2B12# => romdata <= X"818C0000";
    when 16#2B13# => romdata <= X"01000000";
    when 16#2B14# => romdata <= X"01000000";
    when 16#2B15# => romdata <= X"01000000";
    when 16#2B16# => romdata <= X"81C48000";
    when 16#2B17# => romdata <= X"81CCA004";
    when 16#2B18# => romdata <= X"81C3E008";
    when 16#2B19# => romdata <= X"01000000";
    when 16#2B1A# => romdata <= X"81C1E008";
    when 16#2B1B# => romdata <= X"01000000";
    when 16#2B1C# => romdata <= X"A7480000";
    when 16#2B1D# => romdata <= X"8B34E018";
    when 16#2B1E# => romdata <= X"8A096003";
    when 16#2B1F# => romdata <= X"80A16003";
    when 16#2B20# => romdata <= X"12800008";
    when 16#2B21# => romdata <= X"01000000";
    when 16#2B22# => romdata <= X"21100035";
    when 16#2B23# => romdata <= X"A014221C";
    when 16#2B24# => romdata <= X"A2102003";
    when 16#2B25# => romdata <= X"E2240000";
    when 16#2B26# => romdata <= X"8B444000";
    when 16#2B27# => romdata <= X"10800008";
    when 16#2B28# => romdata <= X"21100035";
    when 16#2B29# => romdata <= X"A014221C";
    when 16#2B2A# => romdata <= X"A2102002";
    when 16#2B2B# => romdata <= X"E2240000";
    when 16#2B2C# => romdata <= X"21200000";
    when 16#2B2D# => romdata <= X"E6042024";
    when 16#2B2E# => romdata <= X"8B34E014";
    when 16#2B2F# => romdata <= X"8A09601F";
    when 16#2B30# => romdata <= X"27100035";
    when 16#2B31# => romdata <= X"A614E214";
    when 16#2B32# => romdata <= X"CA24C000";
    when 16#2B33# => romdata <= X"8A016001";
    when 16#2B34# => romdata <= X"27100035";
    when 16#2B35# => romdata <= X"A614E210";
    when 16#2B36# => romdata <= X"CA24C000";
    when 16#2B37# => romdata <= X"27100035";
    when 16#2B38# => romdata <= X"A614E218";
    when 16#2B39# => romdata <= X"8A216002";
    when 16#2B3A# => romdata <= X"CA24C000";
    when 16#2B3B# => romdata <= X"81C3E008";
    when 16#2B3C# => romdata <= X"01000000";
    when 16#2B3D# => romdata <= X"81C3E008";
    when 16#2B3E# => romdata <= X"01000000";
    when 16#2B3F# => romdata <= X"91D02000";
    when 16#2B40# => romdata <= X"01000000";
    when 16#2B41# => romdata <= X"01000000";
    when 16#2B42# => romdata <= X"01000000";
    when 16#2B43# => romdata <= X"81C44000";
    when 16#2B44# => romdata <= X"81CC8000";
    when 16#2B45# => romdata <= X"83480000";
    when 16#2B46# => romdata <= X"83306018";
    when 16#2B47# => romdata <= X"82086003";
    when 16#2B48# => romdata <= X"80A06003";
    when 16#2B49# => romdata <= X"12800006";
    when 16#2B4A# => romdata <= X"01000000";
    when 16#2B4B# => romdata <= X"83444000";
    when 16#2B4C# => romdata <= X"05000008";
    when 16#2B4D# => romdata <= X"82284002";
    when 16#2B4E# => romdata <= X"A3804000";
    when 16#2B4F# => romdata <= X"88100000";
    when 16#2B50# => romdata <= X"0910002A";
    when 16#2B51# => romdata <= X"81C123A4";
    when 16#2B52# => romdata <= X"01000000";
    when 16#2B53# => romdata <= X"9DE3BFA0";
    when 16#2B54# => romdata <= X"21100030";
    when 16#2B55# => romdata <= X"23100030";
    when 16#2B56# => romdata <= X"A01420F8";
    when 16#2B57# => romdata <= X"A21460F8";
    when 16#2B58# => romdata <= X"80A40011";
    when 16#2B59# => romdata <= X"1A80000B";
    when 16#2B5A# => romdata <= X"01000000";
    when 16#2B5B# => romdata <= X"D0040000";
    when 16#2B5C# => romdata <= X"80A22000";
    when 16#2B5D# => romdata <= X"02800004";
    when 16#2B5E# => romdata <= X"A0042004";
    when 16#2B5F# => romdata <= X"9FC20000";
    when 16#2B60# => romdata <= X"01000000";
    when 16#2B61# => romdata <= X"80A40011";
    when 16#2B62# => romdata <= X"2ABFFFFA";
    when 16#2B63# => romdata <= X"D0040000";
    when 16#2B64# => romdata <= X"81C7E008";
    when 16#2B65# => romdata <= X"81E80000";
    when 16#2B66# => romdata <= X"AA27A140";
    when 16#2B67# => romdata <= X"E0256060";
    when 16#2B68# => romdata <= X"E2256064";
    when 16#2B69# => romdata <= X"E4256068";
    when 16#2B6A# => romdata <= X"C2256074";
    when 16#2B6B# => romdata <= X"C43D6078";
    when 16#2B6C# => romdata <= X"C83D6080";
    when 16#2B6D# => romdata <= X"CC3D6088";
    when 16#2B6E# => romdata <= X"85400000";
    when 16#2B6F# => romdata <= X"C425606C";
    when 16#2B70# => romdata <= X"F03D6090";
    when 16#2B71# => romdata <= X"F43D6098";
    when 16#2B72# => romdata <= X"F83D60A0";
    when 16#2B73# => romdata <= X"FC3D60A8";
    when 16#2B74# => romdata <= X"05100035";
    when 16#2B75# => romdata <= X"C600A1F4";
    when 16#2B76# => romdata <= X"C625613C";
    when 16#2B77# => romdata <= X"860560B0";
    when 16#2B78# => romdata <= X"C620A1F4";
    when 16#2B79# => romdata <= X"A8102001";
    when 16#2B7A# => romdata <= X"A92D0010";
    when 16#2B7B# => romdata <= X"808D0013";
    when 16#2B7C# => romdata <= X"02800013";
    when 16#2B7D# => romdata <= X"01000000";
    when 16#2B7E# => romdata <= X"8534E001";
    when 16#2B7F# => romdata <= X"07100035";
    when 16#2B80# => romdata <= X"C600E214";
    when 16#2B81# => romdata <= X"A72CC003";
    when 16#2B82# => romdata <= X"8414C002";
    when 16#2B83# => romdata <= X"8408A0FF";
    when 16#2B84# => romdata <= X"81E00000";
    when 16#2B85# => romdata <= X"8190A000";
    when 16#2B86# => romdata <= X"E03BA000";
    when 16#2B87# => romdata <= X"E43BA008";
    when 16#2B88# => romdata <= X"E83BA010";
    when 16#2B89# => romdata <= X"EC3BA018";
    when 16#2B8A# => romdata <= X"F03BA020";
    when 16#2B8B# => romdata <= X"F43BA028";
    when 16#2B8C# => romdata <= X"F83BA030";
    when 16#2B8D# => romdata <= X"FC3BA038";
    when 16#2B8E# => romdata <= X"81E80000";
    when 16#2B8F# => romdata <= X"81C5A008";
    when 16#2B90# => romdata <= X"9C100015";
    when 16#2B91# => romdata <= X"05100038";
    when 16#2B92# => romdata <= X"8410A23C";
    when 16#2B93# => romdata <= X"C4008000";
    when 16#2B94# => romdata <= X"80A08000";
    when 16#2B95# => romdata <= X"02800004";
    when 16#2B96# => romdata <= X"01000000";
    when 16#2B97# => romdata <= X"9FC08000";
    when 16#2B98# => romdata <= X"9203A0F8";
    when 16#2B99# => romdata <= X"C403A13C";
    when 16#2B9A# => romdata <= X"07100035";
    when 16#2B9B# => romdata <= X"C420E1F4";
    when 16#2B9C# => romdata <= X"818C2000";
    when 16#2B9D# => romdata <= X"82102002";
    when 16#2B9E# => romdata <= X"83284010";
    when 16#2B9F# => romdata <= X"05100035";
    when 16#2BA0# => romdata <= X"C400A210";
    when 16#2BA1# => romdata <= X"85304002";
    when 16#2BA2# => romdata <= X"82104002";
    when 16#2BA3# => romdata <= X"85500000";
    when 16#2BA4# => romdata <= X"80888001";
    when 16#2BA5# => romdata <= X"02800020";
    when 16#2BA6# => romdata <= X"8328A001";
    when 16#2BA7# => romdata <= X"07100035";
    when 16#2BA8# => romdata <= X"C600E214";
    when 16#2BA9# => romdata <= X"85308003";
    when 16#2BAA# => romdata <= X"82104002";
    when 16#2BAB# => romdata <= X"820860FF";
    when 16#2BAC# => romdata <= X"81906000";
    when 16#2BAD# => romdata <= X"C203A06C";
    when 16#2BAE# => romdata <= X"81806000";
    when 16#2BAF# => romdata <= X"F01BA090";
    when 16#2BB0# => romdata <= X"F41BA098";
    when 16#2BB1# => romdata <= X"F81BA0A0";
    when 16#2BB2# => romdata <= X"FC1BA0A8";
    when 16#2BB3# => romdata <= X"C203A074";
    when 16#2BB4# => romdata <= X"C41BA078";
    when 16#2BB5# => romdata <= X"C81BA080";
    when 16#2BB6# => romdata <= X"CC1BA088";
    when 16#2BB7# => romdata <= X"E003A060";
    when 16#2BB8# => romdata <= X"E203A064";
    when 16#2BB9# => romdata <= X"E403A068";
    when 16#2BBA# => romdata <= X"81E80000";
    when 16#2BBB# => romdata <= X"E01BA000";
    when 16#2BBC# => romdata <= X"E41BA008";
    when 16#2BBD# => romdata <= X"E81BA010";
    when 16#2BBE# => romdata <= X"EC1BA018";
    when 16#2BBF# => romdata <= X"F01BA020";
    when 16#2BC0# => romdata <= X"F41BA028";
    when 16#2BC1# => romdata <= X"F81BA030";
    when 16#2BC2# => romdata <= X"FC1BA038";
    when 16#2BC3# => romdata <= X"1080000F";
    when 16#2BC4# => romdata <= X"81E00000";
    when 16#2BC5# => romdata <= X"C203A06C";
    when 16#2BC6# => romdata <= X"81806000";
    when 16#2BC7# => romdata <= X"F01BA090";
    when 16#2BC8# => romdata <= X"F41BA098";
    when 16#2BC9# => romdata <= X"F81BA0A0";
    when 16#2BCA# => romdata <= X"FC1BA0A8";
    when 16#2BCB# => romdata <= X"C203A074";
    when 16#2BCC# => romdata <= X"C41BA078";
    when 16#2BCD# => romdata <= X"C81BA080";
    when 16#2BCE# => romdata <= X"CC1BA088";
    when 16#2BCF# => romdata <= X"E003A060";
    when 16#2BD0# => romdata <= X"E203A064";
    when 16#2BD1# => romdata <= X"E403A068";
    when 16#2BD2# => romdata <= X"818C2000";
    when 16#2BD3# => romdata <= X"01000000";
    when 16#2BD4# => romdata <= X"01000000";
    when 16#2BD5# => romdata <= X"01000000";
    when 16#2BD6# => romdata <= X"81C44000";
    when 16#2BD7# => romdata <= X"81CC8000";
    when 16#2BD8# => romdata <= X"AA27A140";
    when 16#2BD9# => romdata <= X"E0256138";
    when 16#2BDA# => romdata <= X"29000004";
    when 16#2BDB# => romdata <= X"A02C0014";
    when 16#2BDC# => romdata <= X"C2256074";
    when 16#2BDD# => romdata <= X"C43D6078";
    when 16#2BDE# => romdata <= X"C83D6080";
    when 16#2BDF# => romdata <= X"CC3D6088";
    when 16#2BE0# => romdata <= X"85400000";
    when 16#2BE1# => romdata <= X"C425606C";
    when 16#2BE2# => romdata <= X"05100035";
    when 16#2BE3# => romdata <= X"C600A1F4";
    when 16#2BE4# => romdata <= X"C625613C";
    when 16#2BE5# => romdata <= X"860560B0";
    when 16#2BE6# => romdata <= X"C620A1F4";
    when 16#2BE7# => romdata <= X"C020E080";
    when 16#2BE8# => romdata <= X"A8102001";
    when 16#2BE9# => romdata <= X"A92D0010";
    when 16#2BEA# => romdata <= X"808D0013";
    when 16#2BEB# => romdata <= X"02800013";
    when 16#2BEC# => romdata <= X"01000000";
    when 16#2BED# => romdata <= X"8534E001";
    when 16#2BEE# => romdata <= X"07100035";
    when 16#2BEF# => romdata <= X"C600E214";
    when 16#2BF0# => romdata <= X"A72CC003";
    when 16#2BF1# => romdata <= X"8414C002";
    when 16#2BF2# => romdata <= X"8408A0FF";
    when 16#2BF3# => romdata <= X"81E00000";
    when 16#2BF4# => romdata <= X"8190A000";
    when 16#2BF5# => romdata <= X"E03BA000";
    when 16#2BF6# => romdata <= X"E43BA008";
    when 16#2BF7# => romdata <= X"E83BA010";
    when 16#2BF8# => romdata <= X"EC3BA018";
    when 16#2BF9# => romdata <= X"F03BA020";
    when 16#2BFA# => romdata <= X"F43BA028";
    when 16#2BFB# => romdata <= X"F83BA030";
    when 16#2BFC# => romdata <= X"FC3BA038";
    when 16#2BFD# => romdata <= X"81E80000";
    when 16#2BFE# => romdata <= X"81C5A008";
    when 16#2BFF# => romdata <= X"9C100015";
    when 16#2C00# => romdata <= X"05100038";
    when 16#2C01# => romdata <= X"8410A23C";
    when 16#2C02# => romdata <= X"C4008000";
    when 16#2C03# => romdata <= X"80A08000";
    when 16#2C04# => romdata <= X"02800004";
    when 16#2C05# => romdata <= X"01000000";
    when 16#2C06# => romdata <= X"9FC08000";
    when 16#2C07# => romdata <= X"9203A0F8";
    when 16#2C08# => romdata <= X"C403A13C";
    when 16#2C09# => romdata <= X"07100035";
    when 16#2C0A# => romdata <= X"C420E1F4";
    when 16#2C0B# => romdata <= X"07100035";
    when 16#2C0C# => romdata <= X"C600E1F0";
    when 16#2C0D# => romdata <= X"80A08003";
    when 16#2C0E# => romdata <= X"12800008";
    when 16#2C0F# => romdata <= X"01000000";
    when 16#2C10# => romdata <= X"C403A138";
    when 16#2C11# => romdata <= X"07000004";
    when 16#2C12# => romdata <= X"84088003";
    when 16#2C13# => romdata <= X"A02C0003";
    when 16#2C14# => romdata <= X"A0140002";
    when 16#2C15# => romdata <= X"30800006";
    when 16#2C16# => romdata <= X"8403A0B0";
    when 16#2C17# => romdata <= X"80A08003";
    when 16#2C18# => romdata <= X"12800003";
    when 16#2C19# => romdata <= X"07100035";
    when 16#2C1A# => romdata <= X"C020E1F0";
    when 16#2C1B# => romdata <= X"818C2000";
    when 16#2C1C# => romdata <= X"82102002";
    when 16#2C1D# => romdata <= X"83284010";
    when 16#2C1E# => romdata <= X"05100035";
    when 16#2C1F# => romdata <= X"C400A210";
    when 16#2C20# => romdata <= X"85304002";
    when 16#2C21# => romdata <= X"82104002";
    when 16#2C22# => romdata <= X"85500000";
    when 16#2C23# => romdata <= X"80888001";
    when 16#2C24# => romdata <= X"02800019";
    when 16#2C25# => romdata <= X"8328A001";
    when 16#2C26# => romdata <= X"07100035";
    when 16#2C27# => romdata <= X"C600E214";
    when 16#2C28# => romdata <= X"85308003";
    when 16#2C29# => romdata <= X"82104002";
    when 16#2C2A# => romdata <= X"820860FF";
    when 16#2C2B# => romdata <= X"81906000";
    when 16#2C2C# => romdata <= X"C203A06C";
    when 16#2C2D# => romdata <= X"81806000";
    when 16#2C2E# => romdata <= X"C203A074";
    when 16#2C2F# => romdata <= X"C41BA078";
    when 16#2C30# => romdata <= X"C81BA080";
    when 16#2C31# => romdata <= X"CC1BA088";
    when 16#2C32# => romdata <= X"81E80000";
    when 16#2C33# => romdata <= X"E01BA000";
    when 16#2C34# => romdata <= X"E41BA008";
    when 16#2C35# => romdata <= X"E81BA010";
    when 16#2C36# => romdata <= X"EC1BA018";
    when 16#2C37# => romdata <= X"F01BA020";
    when 16#2C38# => romdata <= X"F41BA028";
    when 16#2C39# => romdata <= X"F81BA030";
    when 16#2C3A# => romdata <= X"FC1BA038";
    when 16#2C3B# => romdata <= X"10800008";
    when 16#2C3C# => romdata <= X"81E00000";
    when 16#2C3D# => romdata <= X"C203A06C";
    when 16#2C3E# => romdata <= X"81806000";
    when 16#2C3F# => romdata <= X"C203A074";
    when 16#2C40# => romdata <= X"C41BA078";
    when 16#2C41# => romdata <= X"C81BA080";
    when 16#2C42# => romdata <= X"CC1BA088";
    when 16#2C43# => romdata <= X"818C2000";
    when 16#2C44# => romdata <= X"01000000";
    when 16#2C45# => romdata <= X"01000000";
    when 16#2C46# => romdata <= X"01000000";
    when 16#2C47# => romdata <= X"81C44000";
    when 16#2C48# => romdata <= X"81CC8000";
    when 16#2C49# => romdata <= X"82100008";
    when 16#2C4A# => romdata <= X"9A103800";
    when 16#2C4B# => romdata <= X"96102000";
    when 16#2C4C# => romdata <= X"912AE005";
    when 16#2C4D# => romdata <= X"98034008";
    when 16#2C4E# => romdata <= X"D4034008";
    when 16#2C4F# => romdata <= X"9132A018";
    when 16#2C50# => romdata <= X"80A20001";
    when 16#2C51# => romdata <= X"32800008";
    when 16#2C52# => romdata <= X"9602E001";
    when 16#2C53# => romdata <= X"9132A00C";
    when 16#2C54# => romdata <= X"900A2FFF";
    when 16#2C55# => romdata <= X"80A20009";
    when 16#2C56# => romdata <= X"02800007";
    when 16#2C57# => romdata <= X"9410000C";
    when 16#2C58# => romdata <= X"9602E001";
    when 16#2C59# => romdata <= X"80A2E007";
    when 16#2C5A# => romdata <= X"28BFFFF3";
    when 16#2C5B# => romdata <= X"912AE005";
    when 16#2C5C# => romdata <= X"94102000";
    when 16#2C5D# => romdata <= X"81C3E008";
    when 16#2C5E# => romdata <= X"9010000A";
    when 16#2C5F# => romdata <= X"82100008";
    when 16#2C60# => romdata <= X"98102000";
    when 16#2C61# => romdata <= X"912B2003";
    when 16#2C62# => romdata <= X"9A004008";
    when 16#2C63# => romdata <= X"D6004008";
    when 16#2C64# => romdata <= X"9132E018";
    when 16#2C65# => romdata <= X"80A20009";
    when 16#2C66# => romdata <= X"32800008";
    when 16#2C67# => romdata <= X"98032001";
    when 16#2C68# => romdata <= X"9132E00C";
    when 16#2C69# => romdata <= X"900A2FFF";
    when 16#2C6A# => romdata <= X"80A2000A";
    when 16#2C6B# => romdata <= X"02800007";
    when 16#2C6C# => romdata <= X"9610000D";
    when 16#2C6D# => romdata <= X"98032001";
    when 16#2C6E# => romdata <= X"80A3200F";
    when 16#2C6F# => romdata <= X"28BFFFF3";
    when 16#2C70# => romdata <= X"912B2003";
    when 16#2C71# => romdata <= X"96102000";
    when 16#2C72# => romdata <= X"81C3E008";
    when 16#2C73# => romdata <= X"9010000B";
    when 16#2C74# => romdata <= X"D4022004";
    when 16#2C75# => romdata <= X"173FFC00";
    when 16#2C76# => romdata <= X"920A400B";
    when 16#2C77# => romdata <= X"900A800B";
    when 16#2C78# => romdata <= X"9132200C";
    when 16#2C79# => romdata <= X"92124008";
    when 16#2C7A# => romdata <= X"1100003F";
    when 16#2C7B# => romdata <= X"901223F0";
    when 16#2C7C# => romdata <= X"940A8008";
    when 16#2C7D# => romdata <= X"952AA004";
    when 16#2C7E# => romdata <= X"9412800B";
    when 16#2C7F# => romdata <= X"920A400A";
    when 16#2C80# => romdata <= X"81C3E008";
    when 16#2C81# => romdata <= X"90100009";
    when 16#2C82# => romdata <= X"03100032";
    when 16#2C83# => romdata <= X"81C3E008";
    when 16#2C84# => romdata <= X"D00062C8";
    when 16#2C85# => romdata <= X"9DE3BFA0";
    when 16#2C86# => romdata <= X"21100030";
    when 16#2C87# => romdata <= X"A01420E0";
    when 16#2C88# => romdata <= X"C2043FFC";
    when 16#2C89# => romdata <= X"80A07FFF";
    when 16#2C8A# => romdata <= X"02800008";
    when 16#2C8B# => romdata <= X"A0043FFC";
    when 16#2C8C# => romdata <= X"9FC04000";
    when 16#2C8D# => romdata <= X"A0043FFC";
    when 16#2C8E# => romdata <= X"C2040000";
    when 16#2C8F# => romdata <= X"80A07FFF";
    when 16#2C90# => romdata <= X"12BFFFFC";
    when 16#2C91# => romdata <= X"01000000";
    when 16#2C92# => romdata <= X"81C7E008";
    when 16#2C93# => romdata <= X"81E80000";
    when 16#2C94# => romdata <= X"9DE3BFA0";
    when 16#2C95# => romdata <= X"81C7E008";
    when 16#2C96# => romdata <= X"81E80000";
    when 16#2C98# => romdata <= X"00000010";
    when 16#2C9A# => romdata <= X"017A5200";
    when 16#2C9B# => romdata <= X"047C0F01";
    when 16#2C9C# => romdata <= X"1B0C0E00";
    when 16#2C9D# => romdata <= X"00000010";
    when 16#2C9E# => romdata <= X"00000018";
    when 16#2C9F# => romdata <= X"FFFF5F1C";
    when 16#2CA0# => romdata <= X"00000008";
    when 16#2CA2# => romdata <= X"00000018";
    when 16#2CA4# => romdata <= X"017A5052";
    when 16#2CA5# => romdata <= X"00047C0F";
    when 16#2CA6# => romdata <= X"06004000";
    when 16#2CA7# => romdata <= X"DE781B0C";
    when 16#2CA8# => romdata <= X"0E000000";
    when 16#2CA9# => romdata <= X"00000010";
    when 16#2CAA# => romdata <= X"00000020";
    when 16#2CAB# => romdata <= X"FFFF5EF4";
    when 16#2CAC# => romdata <= X"0000000C";
    when 16#2CAE# => romdata <= X"00000010";
    when 16#2CAF# => romdata <= X"00000034";
    when 16#2CB0# => romdata <= X"FFFF5EEC";
    when 16#2CB1# => romdata <= X"0000000C";
    when 16#2CB3# => romdata <= X"00000018";
    when 16#2CB4# => romdata <= X"00000048";
    when 16#2CB5# => romdata <= X"FFFF5EE4";
    when 16#2CB6# => romdata <= X"0000008C";
    when 16#2CB7# => romdata <= X"00410D1E";
    when 16#2CB8# => romdata <= X"2D4D090F";
    when 16#2CB9# => romdata <= X"1F000000";
    when 16#2CBA# => romdata <= X"00000018";
    when 16#2CBB# => romdata <= X"00000064";
    when 16#2CBC# => romdata <= X"FFFF5F54";
    when 16#2CBD# => romdata <= X"000000B8";
    when 16#2CBE# => romdata <= X"00410D1E";
    when 16#2CBF# => romdata <= X"2D41090F";
    when 16#2CC0# => romdata <= X"1F000000";
    when 16#2CC1# => romdata <= X"00000010";
    when 16#2CC2# => romdata <= X"00000080";
    when 16#2CC3# => romdata <= X"FFFF5FF0";
    when 16#2CC4# => romdata <= X"00000020";
    when 16#2CC6# => romdata <= X"00000010";
    when 16#2CC7# => romdata <= X"00000094";
    when 16#2CC8# => romdata <= X"FFFF5FFC";
    when 16#2CC9# => romdata <= X"00000014";
    when 16#2CCB# => romdata <= X"00000010";
    when 16#2CCC# => romdata <= X"000000A8";
    when 16#2CCD# => romdata <= X"FFFF5FFC";
    when 16#2CCE# => romdata <= X"00000028";
    when 16#2CD0# => romdata <= X"00000010";
    when 16#2CD1# => romdata <= X"000000BC";
    when 16#2CD2# => romdata <= X"FFFF6010";
    when 16#2CD3# => romdata <= X"0000006C";
    when 16#2CD5# => romdata <= X"00000018";
    when 16#2CD6# => romdata <= X"000000D0";
    when 16#2CD7# => romdata <= X"FFFF6068";
    when 16#2CD8# => romdata <= X"0000004C";
    when 16#2CD9# => romdata <= X"00410D1E";
    when 16#2CDA# => romdata <= X"2D4A090F";
    when 16#2CDB# => romdata <= X"1F000000";
    when 16#2CDC# => romdata <= X"00000010";
    when 16#2CDD# => romdata <= X"000000EC";
    when 16#2CDE# => romdata <= X"FFFF6098";
    when 16#2CDF# => romdata <= X"0000000C";
    when 16#2CE1# => romdata <= X"00000010";
    when 16#2CE2# => romdata <= X"00000100";
    when 16#2CE3# => romdata <= X"FFFF6090";
    when 16#2CE4# => romdata <= X"0000000C";
    when 16#2CE6# => romdata <= X"00000010";
    when 16#2CE7# => romdata <= X"00000114";
    when 16#2CE8# => romdata <= X"FFFF6088";
    when 16#2CE9# => romdata <= X"00000010";
    when 16#2CEB# => romdata <= X"00000010";
    when 16#2CEC# => romdata <= X"00000128";
    when 16#2CED# => romdata <= X"FFFF6084";
    when 16#2CEE# => romdata <= X"0000002C";
    when 16#2CF0# => romdata <= X"00000010";
    when 16#2CF1# => romdata <= X"0000013C";
    when 16#2CF2# => romdata <= X"FFFF609C";
    when 16#2CF3# => romdata <= X"0000002C";
    when 16#2CF5# => romdata <= X"00000010";
    when 16#2CF6# => romdata <= X"00000150";
    when 16#2CF7# => romdata <= X"FFFF60E0";
    when 16#2CF8# => romdata <= X"00000048";
    when 16#2CFA# => romdata <= X"00000018";
    when 16#2CFB# => romdata <= X"00000164";
    when 16#2CFC# => romdata <= X"FFFF6114";
    when 16#2CFD# => romdata <= X"000002E0";
    when 16#2CFE# => romdata <= X"00410D1E";
    when 16#2CFF# => romdata <= X"2D4B090F";
    when 16#2D00# => romdata <= X"1F000000";
    when 16#2D01# => romdata <= X"00000018";
    when 16#2D02# => romdata <= X"00000180";
    when 16#2D03# => romdata <= X"FFFF63D8";
    when 16#2D04# => romdata <= X"00000290";
    when 16#2D05# => romdata <= X"00410D1E";
    when 16#2D06# => romdata <= X"2D42090F";
    when 16#2D07# => romdata <= X"1F000000";
    when 16#2D08# => romdata <= X"00000010";
    when 16#2D09# => romdata <= X"0000019C";
    when 16#2D0A# => romdata <= X"FFFF666C";
    when 16#2D0B# => romdata <= X"00000008";
    when 16#2D0D# => romdata <= X"00000010";
    when 16#2D0E# => romdata <= X"000001B0";
    when 16#2D0F# => romdata <= X"FFFF6660";
    when 16#2D10# => romdata <= X"0000003C";
    when 16#2D12# => romdata <= X"00000010";
    when 16#2D13# => romdata <= X"000001C4";
    when 16#2D14# => romdata <= X"FFFF6688";
    when 16#2D15# => romdata <= X"00000050";
    when 16#2D17# => romdata <= X"00000018";
    when 16#2D18# => romdata <= X"000001D8";
    when 16#2D19# => romdata <= X"FFFF66C4";
    when 16#2D1A# => romdata <= X"00000028";
    when 16#2D1B# => romdata <= X"00410D1E";
    when 16#2D1C# => romdata <= X"2D45090F";
    when 16#2D1D# => romdata <= X"1F000000";
    when 16#2D1E# => romdata <= X"00000018";
    when 16#2D1F# => romdata <= X"000001F4";
    when 16#2D20# => romdata <= X"FFFF66D0";
    when 16#2D21# => romdata <= X"00000084";
    when 16#2D22# => romdata <= X"00410D1E";
    when 16#2D23# => romdata <= X"2D41090F";
    when 16#2D24# => romdata <= X"1F000000";
    when 16#2D25# => romdata <= X"00000018";
    when 16#2D26# => romdata <= X"00000210";
    when 16#2D27# => romdata <= X"FFFF6738";
    when 16#2D28# => romdata <= X"00000064";
    when 16#2D29# => romdata <= X"00410D1E";
    when 16#2D2A# => romdata <= X"2D41090F";
    when 16#2D2B# => romdata <= X"1F000000";
    when 16#2D2C# => romdata <= X"00000018";
    when 16#2D2D# => romdata <= X"0000022C";
    when 16#2D2E# => romdata <= X"FFFF6780";
    when 16#2D2F# => romdata <= X"000003C8";
    when 16#2D30# => romdata <= X"00410D1E";
    when 16#2D31# => romdata <= X"2D47090F";
    when 16#2D32# => romdata <= X"1F000000";
    when 16#2D33# => romdata <= X"00000014";
    when 16#2D34# => romdata <= X"00000248";
    when 16#2D35# => romdata <= X"FFFF6B2C";
    when 16#2D36# => romdata <= X"0000009C";
    when 16#2D37# => romdata <= X"00410D1E";
    when 16#2D38# => romdata <= X"2D090F1F";
    when 16#2D39# => romdata <= X"00000014";
    when 16#2D3A# => romdata <= X"00000260";
    when 16#2D3B# => romdata <= X"FFFF6BB0";
    when 16#2D3C# => romdata <= X"000000A4";
    when 16#2D3D# => romdata <= X"00410D1E";
    when 16#2D3E# => romdata <= X"2D090F1F";
    when 16#2D3F# => romdata <= X"00000018";
    when 16#2D40# => romdata <= X"00000278";
    when 16#2D41# => romdata <= X"FFFF6C3C";
    when 16#2D42# => romdata <= X"0000010C";
    when 16#2D43# => romdata <= X"00410D1E";
    when 16#2D44# => romdata <= X"2D43090F";
    when 16#2D45# => romdata <= X"1F000000";
    when 16#2D46# => romdata <= X"00000018";
    when 16#2D47# => romdata <= X"00000294";
    when 16#2D48# => romdata <= X"FFFF6D2C";
    when 16#2D49# => romdata <= X"0000014C";
    when 16#2D4A# => romdata <= X"00410D1E";
    when 16#2D4B# => romdata <= X"2D4E090F";
    when 16#2D4C# => romdata <= X"1F000000";
    when 16#2D4D# => romdata <= X"00000010";
    when 16#2D4E# => romdata <= X"000002B0";
    when 16#2D4F# => romdata <= X"FFFF6E5C";
    when 16#2D50# => romdata <= X"00000008";
    when 16#2D52# => romdata <= X"00000010";
    when 16#2D53# => romdata <= X"000002C4";
    when 16#2D54# => romdata <= X"FFFF6E50";
    when 16#2D55# => romdata <= X"00000008";
    when 16#2D57# => romdata <= X"00000010";
    when 16#2D58# => romdata <= X"000002D8";
    when 16#2D59# => romdata <= X"FFFF6E44";
    when 16#2D5A# => romdata <= X"00000008";
    when 16#2D5C# => romdata <= X"00000010";
    when 16#2D5D# => romdata <= X"000002EC";
    when 16#2D5E# => romdata <= X"FFFF6E38";
    when 16#2D5F# => romdata <= X"00000008";
    when 16#2D61# => romdata <= X"00000010";
    when 16#2D62# => romdata <= X"00000300";
    when 16#2D63# => romdata <= X"FFFF6E2C";
    when 16#2D64# => romdata <= X"00000040";
    when 16#2D66# => romdata <= X"00000010";
    when 16#2D67# => romdata <= X"00000314";
    when 16#2D68# => romdata <= X"FFFF6E58";
    when 16#2D69# => romdata <= X"00000028";
    when 16#2D6B# => romdata <= X"00000018";
    when 16#2D6C# => romdata <= X"00000328";
    when 16#2D6D# => romdata <= X"FFFF6E6C";
    when 16#2D6E# => romdata <= X"000000DC";
    when 16#2D6F# => romdata <= X"00410D1E";
    when 16#2D70# => romdata <= X"2D66090F";
    when 16#2D71# => romdata <= X"1F000000";
    when 16#2D72# => romdata <= X"00000018";
    when 16#2D73# => romdata <= X"00000344";
    when 16#2D74# => romdata <= X"FFFF6F2C";
    when 16#2D75# => romdata <= X"0000002C";
    when 16#2D76# => romdata <= X"00410D1E";
    when 16#2D77# => romdata <= X"2D44090F";
    when 16#2D78# => romdata <= X"1F000000";
    when 16#2D79# => romdata <= X"00000018";
    when 16#2D7A# => romdata <= X"00000360";
    when 16#2D7B# => romdata <= X"FFFF6F3C";
    when 16#2D7C# => romdata <= X"00000048";
    when 16#2D7D# => romdata <= X"00410D1E";
    when 16#2D7E# => romdata <= X"2D41090F";
    when 16#2D7F# => romdata <= X"1F000000";
    when 16#2D80# => romdata <= X"00000010";
    when 16#2D81# => romdata <= X"000003A4";
    when 16#2D82# => romdata <= X"FFFF6F68";
    when 16#2D83# => romdata <= X"00000020";
    when 16#2D85# => romdata <= X"00000010";
    when 16#2D86# => romdata <= X"000003B8";
    when 16#2D87# => romdata <= X"FFFF6F74";
    when 16#2D88# => romdata <= X"00000024";
    when 16#2D8A# => romdata <= X"00000010";
    when 16#2D8B# => romdata <= X"000003CC";
    when 16#2D8C# => romdata <= X"FFFF6F84";
    when 16#2D8D# => romdata <= X"000000E8";
    when 16#2D8F# => romdata <= X"00000018";
    when 16#2D90# => romdata <= X"000003E0";
    when 16#2D91# => romdata <= X"FFFF7058";
    when 16#2D92# => romdata <= X"00000050";
    when 16#2D93# => romdata <= X"00410D1E";
    when 16#2D94# => romdata <= X"2D4D090F";
    when 16#2D95# => romdata <= X"1F000000";
    when 16#2D96# => romdata <= X"00000018";
    when 16#2D97# => romdata <= X"000003FC";
    when 16#2D98# => romdata <= X"FFFF708C";
    when 16#2D99# => romdata <= X"00000054";
    when 16#2D9A# => romdata <= X"00410D1E";
    when 16#2D9B# => romdata <= X"2D4E090F";
    when 16#2D9C# => romdata <= X"1F000000";
    when 16#2D9D# => romdata <= X"00000018";
    when 16#2D9E# => romdata <= X"00000418";
    when 16#2D9F# => romdata <= X"FFFF70C4";
    when 16#2DA0# => romdata <= X"0000012C";
    when 16#2DA1# => romdata <= X"00410D1E";
    when 16#2DA2# => romdata <= X"2D41090F";
    when 16#2DA3# => romdata <= X"1F000000";
    when 16#2DA4# => romdata <= X"00000010";
    when 16#2DA5# => romdata <= X"00000434";
    when 16#2DA6# => romdata <= X"FFFF71D4";
    when 16#2DA7# => romdata <= X"0000001C";
    when 16#2DA9# => romdata <= X"00000010";
    when 16#2DAA# => romdata <= X"00000448";
    when 16#2DAB# => romdata <= X"FFFF71DC";
    when 16#2DAC# => romdata <= X"0000001C";
    when 16#2DAE# => romdata <= X"00000018";
    when 16#2DAF# => romdata <= X"0000045C";
    when 16#2DB0# => romdata <= X"FFFF71E4";
    when 16#2DB1# => romdata <= X"000006D8";
    when 16#2DB2# => romdata <= X"00410D1E";
    when 16#2DB3# => romdata <= X"2D4C090F";
    when 16#2DB4# => romdata <= X"1F000000";
    when 16#2DB5# => romdata <= X"00000010";
    when 16#2DB6# => romdata <= X"00000478";
    when 16#2DB7# => romdata <= X"FFFF78A0";
    when 16#2DB8# => romdata <= X"00000018";
    when 16#2DBA# => romdata <= X"00000010";
    when 16#2DBB# => romdata <= X"0000048C";
    when 16#2DBC# => romdata <= X"FFFF78A4";
    when 16#2DBD# => romdata <= X"00000018";
    when 16#2DBF# => romdata <= X"00000018";
    when 16#2DC0# => romdata <= X"000004A0";
    when 16#2DC1# => romdata <= X"FFFF78A8";
    when 16#2DC2# => romdata <= X"00000040";
    when 16#2DC3# => romdata <= X"00410D1E";
    when 16#2DC4# => romdata <= X"2D42090F";
    when 16#2DC5# => romdata <= X"1F000000";
    when 16#2DC6# => romdata <= X"00000018";
    when 16#2DC7# => romdata <= X"000004BC";
    when 16#2DC8# => romdata <= X"FFFF7A30";
    when 16#2DC9# => romdata <= X"00000038";
    when 16#2DCA# => romdata <= X"00410D1E";
    when 16#2DCB# => romdata <= X"2D47090F";
    when 16#2DCC# => romdata <= X"1F000000";
    when 16#2DCD# => romdata <= X"00000014";
    when 16#2DCE# => romdata <= X"000004D8";
    when 16#2DCF# => romdata <= X"FFFF7A4C";
    when 16#2DD0# => romdata <= X"00001D54";
    when 16#2DD1# => romdata <= X"00410D1E";
    when 16#2DD2# => romdata <= X"2D090F1F";
    when 16#2DD3# => romdata <= X"00000010";
    when 16#2DD4# => romdata <= X"000004F0";
    when 16#2DD5# => romdata <= X"FFFF9788";
    when 16#2DD6# => romdata <= X"0000002C";
    when 16#2DD8# => romdata <= X"00000018";
    when 16#2DD9# => romdata <= X"00000504";
    when 16#2DDA# => romdata <= X"FFFF97A0";
    when 16#2DDB# => romdata <= X"00000060";
    when 16#2DDC# => romdata <= X"00410D1E";
    when 16#2DDD# => romdata <= X"2D46090F";
    when 16#2DDE# => romdata <= X"1F000000";
    when 16#2DDF# => romdata <= X"00000010";
    when 16#2DE0# => romdata <= X"00000520";
    when 16#2DE1# => romdata <= X"FFFF97E4";
    when 16#2DE2# => romdata <= X"0000002C";
    when 16#2DE4# => romdata <= X"00000018";
    when 16#2DE5# => romdata <= X"00000534";
    when 16#2DE6# => romdata <= X"FFFF97FC";
    when 16#2DE7# => romdata <= X"00000138";
    when 16#2DE8# => romdata <= X"00410D1E";
    when 16#2DE9# => romdata <= X"2D4D090F";
    when 16#2DEA# => romdata <= X"1F000000";
    when 16#2DEB# => romdata <= X"00000010";
    when 16#2DEC# => romdata <= X"00000550";
    when 16#2DED# => romdata <= X"FFFF9918";
    when 16#2DEE# => romdata <= X"00000034";
    when 16#2DF0# => romdata <= X"00000018";
    when 16#2DF1# => romdata <= X"00000564";
    when 16#2DF2# => romdata <= X"FFFF9938";
    when 16#2DF3# => romdata <= X"000003F4";
    when 16#2DF4# => romdata <= X"00410D1E";
    when 16#2DF5# => romdata <= X"2D41090F";
    when 16#2DF6# => romdata <= X"1F000000";
    when 16#2DF7# => romdata <= X"00000018";
    when 16#2DF8# => romdata <= X"00000580";
    when 16#2DF9# => romdata <= X"FFFF9D10";
    when 16#2DFA# => romdata <= X"00000134";
    when 16#2DFB# => romdata <= X"00410D1E";
    when 16#2DFC# => romdata <= X"2D49090F";
    when 16#2DFD# => romdata <= X"1F000000";
    when 16#2DFE# => romdata <= X"00000018";
    when 16#2DFF# => romdata <= X"0000059C";
    when 16#2E00# => romdata <= X"FFFF9E28";
    when 16#2E01# => romdata <= X"00000218";
    when 16#2E02# => romdata <= X"00410D1E";
    when 16#2E03# => romdata <= X"2D4E090F";
    when 16#2E04# => romdata <= X"1F000000";
    when 16#2E05# => romdata <= X"00000018";
    when 16#2E06# => romdata <= X"000005B8";
    when 16#2E07# => romdata <= X"FFFFA024";
    when 16#2E08# => romdata <= X"00001304";
    when 16#2E09# => romdata <= X"00410D1E";
    when 16#2E0A# => romdata <= X"2D51090F";
    when 16#2E0B# => romdata <= X"1F000000";
    when 16#2E0C# => romdata <= X"00000018";
    when 16#2E0D# => romdata <= X"000005D4";
    when 16#2E0E# => romdata <= X"FFFFB30C";
    when 16#2E0F# => romdata <= X"0000015C";
    when 16#2E10# => romdata <= X"00410D1E";
    when 16#2E11# => romdata <= X"2D47090F";
    when 16#2E12# => romdata <= X"1F000000";
    when 16#2E13# => romdata <= X"00000010";
    when 16#2E14# => romdata <= X"000005F0";
    when 16#2E15# => romdata <= X"FFFFB44C";
    when 16#2E16# => romdata <= X"00000018";
    when 16#2E18# => romdata <= X"00000010";
    when 16#2E19# => romdata <= X"00000604";
    when 16#2E1A# => romdata <= X"FFFFB450";
    when 16#2E1B# => romdata <= X"00000018";
    when 16#2E1D# => romdata <= X"00000018";
    when 16#2E1E# => romdata <= X"00000618";
    when 16#2E1F# => romdata <= X"FFFFB454";
    when 16#2E20# => romdata <= X"00000024";
    when 16#2E21# => romdata <= X"00410D1E";
    when 16#2E22# => romdata <= X"2D44090F";
    when 16#2E23# => romdata <= X"1F000000";
    when 16#2E24# => romdata <= X"00000010";
    when 16#2E25# => romdata <= X"00000634";
    when 16#2E26# => romdata <= X"FFFFB45C";
    when 16#2E27# => romdata <= X"00000018";
    when 16#2E29# => romdata <= X"00000018";
    when 16#2E2A# => romdata <= X"00000648";
    when 16#2E2B# => romdata <= X"FFFFB460";
    when 16#2E2C# => romdata <= X"00000024";
    when 16#2E2D# => romdata <= X"00410D1E";
    when 16#2E2E# => romdata <= X"2D43090F";
    when 16#2E2F# => romdata <= X"1F000000";
    when 16#2E30# => romdata <= X"00000018";
    when 16#2E31# => romdata <= X"00000664";
    when 16#2E32# => romdata <= X"FFFFB468";
    when 16#2E33# => romdata <= X"00000024";
    when 16#2E34# => romdata <= X"00410D1E";
    when 16#2E35# => romdata <= X"2D44090F";
    when 16#2E36# => romdata <= X"1F000000";
    when 16#2E37# => romdata <= X"00000010";
    when 16#2E38# => romdata <= X"00000680";
    when 16#2E39# => romdata <= X"FFFFB470";
    when 16#2E3A# => romdata <= X"00000018";
    when 16#2E3C# => romdata <= X"00000014";
    when 16#2E3D# => romdata <= X"00000694";
    when 16#2E3E# => romdata <= X"FFFFB474";
    when 16#2E3F# => romdata <= X"00000020";
    when 16#2E40# => romdata <= X"00410D1E";
    when 16#2E41# => romdata <= X"2D090F1F";
    when 16#2E42# => romdata <= X"00000018";
    when 16#2E43# => romdata <= X"000006AC";
    when 16#2E44# => romdata <= X"FFFFB47C";
    when 16#2E45# => romdata <= X"0000008C";
    when 16#2E46# => romdata <= X"00410D1E";
    when 16#2E47# => romdata <= X"2D56090F";
    when 16#2E48# => romdata <= X"1F000000";
    when 16#2E49# => romdata <= X"00000018";
    when 16#2E4A# => romdata <= X"000006C8";
    when 16#2E4B# => romdata <= X"FFFFB4EC";
    when 16#2E4C# => romdata <= X"0000006C";
    when 16#2E4D# => romdata <= X"00410D1E";
    when 16#2E4E# => romdata <= X"2D4D090F";
    when 16#2E4F# => romdata <= X"1F000000";
    when 16#2E50# => romdata <= X"00000018";
    when 16#2E51# => romdata <= X"000006E4";
    when 16#2E52# => romdata <= X"FFFFB53C";
    when 16#2E53# => romdata <= X"00000050";
    when 16#2E54# => romdata <= X"00410D1E";
    when 16#2E55# => romdata <= X"2D46090F";
    when 16#2E56# => romdata <= X"1F000000";
    when 16#2E57# => romdata <= X"00000014";
    when 16#2E58# => romdata <= X"00000700";
    when 16#2E59# => romdata <= X"FFFFB570";
    when 16#2E5A# => romdata <= X"0000011C";
    when 16#2E5B# => romdata <= X"00410D1E";
    when 16#2E5C# => romdata <= X"2D090F1F";
    when 16#2E5D# => romdata <= X"00000014";
    when 16#2E5E# => romdata <= X"00000718";
    when 16#2E5F# => romdata <= X"FFFFB674";
    when 16#2E60# => romdata <= X"000000EC";
    when 16#2E61# => romdata <= X"00410D1E";
    when 16#2E62# => romdata <= X"2D090F1F";
    when 16#2E63# => romdata <= X"00000018";
    when 16#2E64# => romdata <= X"00000730";
    when 16#2E65# => romdata <= X"FFFFB748";
    when 16#2E66# => romdata <= X"0000029C";
    when 16#2E67# => romdata <= X"00410D1E";
    when 16#2E68# => romdata <= X"2D43090F";
    when 16#2E69# => romdata <= X"1F000000";
    when 16#2E6A# => romdata <= X"00000018";
    when 16#2E6B# => romdata <= X"0000074C";
    when 16#2E6C# => romdata <= X"FFFFB9C8";
    when 16#2E6D# => romdata <= X"00000420";
    when 16#2E6E# => romdata <= X"00410D1E";
    when 16#2E6F# => romdata <= X"2D59090F";
    when 16#2E70# => romdata <= X"1F000000";
    when 16#2E71# => romdata <= X"00000014";
    when 16#2E72# => romdata <= X"00000768";
    when 16#2E73# => romdata <= X"FFFFBDCC";
    when 16#2E74# => romdata <= X"000000E4";
    when 16#2E75# => romdata <= X"00410D1E";
    when 16#2E76# => romdata <= X"2D090F1F";
    when 16#2E77# => romdata <= X"00000014";
    when 16#2E78# => romdata <= X"00000780";
    when 16#2E79# => romdata <= X"FFFFBE98";
    when 16#2E7A# => romdata <= X"000000E0";
    when 16#2E7B# => romdata <= X"00410D1E";
    when 16#2E7C# => romdata <= X"2D090F1F";
    when 16#2E7D# => romdata <= X"00000010";
    when 16#2E7E# => romdata <= X"00000798";
    when 16#2E7F# => romdata <= X"FFFFBF60";
    when 16#2E80# => romdata <= X"0000000C";
    when 16#2E82# => romdata <= X"00000010";
    when 16#2E83# => romdata <= X"000007AC";
    when 16#2E84# => romdata <= X"FFFFBF58";
    when 16#2E85# => romdata <= X"0000000C";
    when 16#2E87# => romdata <= X"00000010";
    when 16#2E88# => romdata <= X"000007C0";
    when 16#2E89# => romdata <= X"FFFFBF50";
    when 16#2E8A# => romdata <= X"0000000C";
    when 16#2E8C# => romdata <= X"00000018";
    when 16#2E8D# => romdata <= X"000007D4";
    when 16#2E8E# => romdata <= X"FFFFBF48";
    when 16#2E8F# => romdata <= X"00000068";
    when 16#2E90# => romdata <= X"00410D1E";
    when 16#2E91# => romdata <= X"2D47090F";
    when 16#2E92# => romdata <= X"1F000000";
    when 16#2E93# => romdata <= X"00000010";
    when 16#2E94# => romdata <= X"000007F0";
    when 16#2E95# => romdata <= X"FFFFBF94";
    when 16#2E96# => romdata <= X"00000024";
    when 16#2E98# => romdata <= X"00000018";
    when 16#2E99# => romdata <= X"00000804";
    when 16#2E9A# => romdata <= X"FFFFBFA4";
    when 16#2E9B# => romdata <= X"00000160";
    when 16#2E9C# => romdata <= X"00410D1E";
    when 16#2E9D# => romdata <= X"2D49090F";
    when 16#2E9E# => romdata <= X"1F000000";
    when 16#2E9F# => romdata <= X"00000018";
    when 16#2EA0# => romdata <= X"00000820";
    when 16#2EA1# => romdata <= X"FFFFC0E8";
    when 16#2EA2# => romdata <= X"000000F0";
    when 16#2EA3# => romdata <= X"00410D1E";
    when 16#2EA4# => romdata <= X"2D5B090F";
    when 16#2EA5# => romdata <= X"1F000000";
    when 16#2EA6# => romdata <= X"00000018";
    when 16#2EA7# => romdata <= X"0000083C";
    when 16#2EA8# => romdata <= X"FFFFC1BC";
    when 16#2EA9# => romdata <= X"000000FC";
    when 16#2EAA# => romdata <= X"00410D1E";
    when 16#2EAB# => romdata <= X"2D54090F";
    when 16#2EAC# => romdata <= X"1F000000";
    when 16#2EAD# => romdata <= X"00000018";
    when 16#2EAE# => romdata <= X"00000858";
    when 16#2EAF# => romdata <= X"FFFFC29C";
    when 16#2EB0# => romdata <= X"00000150";
    when 16#2EB1# => romdata <= X"00410D1E";
    when 16#2EB2# => romdata <= X"2D56090F";
    when 16#2EB3# => romdata <= X"1F000000";
    when 16#2EB4# => romdata <= X"00000018";
    when 16#2EB5# => romdata <= X"00000874";
    when 16#2EB6# => romdata <= X"FFFFC3D0";
    when 16#2EB7# => romdata <= X"000000DC";
    when 16#2EB8# => romdata <= X"00410D1E";
    when 16#2EB9# => romdata <= X"2D76090F";
    when 16#2EBA# => romdata <= X"1F000000";
    when 16#2EBB# => romdata <= X"00000010";
    when 16#2EBC# => romdata <= X"00000890";
    when 16#2EBD# => romdata <= X"FFFFC490";
    when 16#2EBE# => romdata <= X"0000002C";
    when 16#2EC0# => romdata <= X"00000010";
    when 16#2EC1# => romdata <= X"000008A4";
    when 16#2EC2# => romdata <= X"FFFFC4A8";
    when 16#2EC3# => romdata <= X"00000084";
    when 16#2EC5# => romdata <= X"00000010";
    when 16#2EC6# => romdata <= X"000008B8";
    when 16#2EC7# => romdata <= X"FFFFC518";
    when 16#2EC8# => romdata <= X"000000E4";
    when 16#2ECA# => romdata <= X"00000018";
    when 16#2ECB# => romdata <= X"000008CC";
    when 16#2ECC# => romdata <= X"FFFFC5E8";
    when 16#2ECD# => romdata <= X"00000074";
    when 16#2ECE# => romdata <= X"00410D1E";
    when 16#2ECF# => romdata <= X"2D57090F";
    when 16#2ED0# => romdata <= X"1F000000";
    when 16#2ED1# => romdata <= X"00000010";
    when 16#2ED2# => romdata <= X"000008E8";
    when 16#2ED3# => romdata <= X"FFFFC640";
    when 16#2ED4# => romdata <= X"0000009C";
    when 16#2ED5# => romdata <= X"00450E68";
    when 16#2ED6# => romdata <= X"00000018";
    when 16#2ED7# => romdata <= X"000008FC";
    when 16#2ED8# => romdata <= X"FFFFC6C8";
    when 16#2ED9# => romdata <= X"00000110";
    when 16#2EDA# => romdata <= X"00410D1E";
    when 16#2EDB# => romdata <= X"2D44090F";
    when 16#2EDC# => romdata <= X"1F000000";
    when 16#2EDD# => romdata <= X"00000018";
    when 16#2EDE# => romdata <= X"00000918";
    when 16#2EDF# => romdata <= X"FFFFC7BC";
    when 16#2EE0# => romdata <= X"000000AC";
    when 16#2EE1# => romdata <= X"00410D1E";
    when 16#2EE2# => romdata <= X"2D41090F";
    when 16#2EE3# => romdata <= X"1F000000";
    when 16#2EE4# => romdata <= X"00000010";
    when 16#2EE5# => romdata <= X"00000934";
    when 16#2EE6# => romdata <= X"FFFFC84C";
    when 16#2EE7# => romdata <= X"00000040";
    when 16#2EE9# => romdata <= X"00000018";
    when 16#2EEA# => romdata <= X"00000948";
    when 16#2EEB# => romdata <= X"FFFFC878";
    when 16#2EEC# => romdata <= X"000000A8";
    when 16#2EED# => romdata <= X"00410D1E";
    when 16#2EEE# => romdata <= X"2D4F090F";
    when 16#2EEF# => romdata <= X"1F000000";
    when 16#2EF0# => romdata <= X"00000018";
    when 16#2EF1# => romdata <= X"00000964";
    when 16#2EF2# => romdata <= X"FFFFC904";
    when 16#2EF3# => romdata <= X"00000130";
    when 16#2EF4# => romdata <= X"00410D1E";
    when 16#2EF5# => romdata <= X"2D43090F";
    when 16#2EF6# => romdata <= X"1F000000";
    when 16#2EF7# => romdata <= X"00000018";
    when 16#2EF8# => romdata <= X"00000980";
    when 16#2EF9# => romdata <= X"FFFFCA18";
    when 16#2EFA# => romdata <= X"000001B4";
    when 16#2EFB# => romdata <= X"00410D1E";
    when 16#2EFC# => romdata <= X"2D4A090F";
    when 16#2EFD# => romdata <= X"1F000000";
    when 16#2EFE# => romdata <= X"00000018";
    when 16#2EFF# => romdata <= X"0000099C";
    when 16#2F00# => romdata <= X"FFFFCBB0";
    when 16#2F01# => romdata <= X"00000134";
    when 16#2F02# => romdata <= X"00410D1E";
    when 16#2F03# => romdata <= X"2D4D090F";
    when 16#2F04# => romdata <= X"1F000000";
    when 16#2F05# => romdata <= X"00000018";
    when 16#2F06# => romdata <= X"000009B8";
    when 16#2F07# => romdata <= X"FFFFCCC8";
    when 16#2F08# => romdata <= X"00000220";
    when 16#2F09# => romdata <= X"00410D1E";
    when 16#2F0A# => romdata <= X"2D4E090F";
    when 16#2F0B# => romdata <= X"1F000000";
    when 16#2F0C# => romdata <= X"00000018";
    when 16#2F0D# => romdata <= X"000009D4";
    when 16#2F0E# => romdata <= X"FFFFCECC";
    when 16#2F0F# => romdata <= X"00000024";
    when 16#2F10# => romdata <= X"00410D1E";
    when 16#2F11# => romdata <= X"2D41090F";
    when 16#2F12# => romdata <= X"1F000000";
    when 16#2F13# => romdata <= X"00000018";
    when 16#2F14# => romdata <= X"000009F0";
    when 16#2F15# => romdata <= X"FFFFCED4";
    when 16#2F16# => romdata <= X"000000E8";
    when 16#2F17# => romdata <= X"00410D1E";
    when 16#2F18# => romdata <= X"2D47090F";
    when 16#2F19# => romdata <= X"1F000000";
    when 16#2F1A# => romdata <= X"00000018";
    when 16#2F1B# => romdata <= X"00000A0C";
    when 16#2F1C# => romdata <= X"FFFFCFA0";
    when 16#2F1D# => romdata <= X"00000114";
    when 16#2F1E# => romdata <= X"00410D1E";
    when 16#2F1F# => romdata <= X"2D47090F";
    when 16#2F20# => romdata <= X"1F000000";
    when 16#2F21# => romdata <= X"00000018";
    when 16#2F22# => romdata <= X"00000A28";
    when 16#2F23# => romdata <= X"FFFFD098";
    when 16#2F24# => romdata <= X"000000D0";
    when 16#2F25# => romdata <= X"00410D1E";
    when 16#2F26# => romdata <= X"2D41090F";
    when 16#2F27# => romdata <= X"1F000000";
    when 16#2F28# => romdata <= X"00000018";
    when 16#2F29# => romdata <= X"00000A44";
    when 16#2F2A# => romdata <= X"FFFFD14C";
    when 16#2F2B# => romdata <= X"000004F8";
    when 16#2F2C# => romdata <= X"00410D1E";
    when 16#2F2D# => romdata <= X"2D43090F";
    when 16#2F2E# => romdata <= X"1F000000";
    when 16#2F2F# => romdata <= X"00000018";
    when 16#2F30# => romdata <= X"00000A60";
    when 16#2F31# => romdata <= X"FFFFD628";
    when 16#2F32# => romdata <= X"0000008C";
    when 16#2F33# => romdata <= X"00410D1E";
    when 16#2F34# => romdata <= X"2D4F090F";
    when 16#2F35# => romdata <= X"1F000000";
    when 16#2F36# => romdata <= X"00000018";
    when 16#2F37# => romdata <= X"00000A7C";
    when 16#2F38# => romdata <= X"FFFFD698";
    when 16#2F39# => romdata <= X"00000028";
    when 16#2F3A# => romdata <= X"00410D1E";
    when 16#2F3B# => romdata <= X"2D44090F";
    when 16#2F3C# => romdata <= X"1F000000";
    when 16#2F3D# => romdata <= X"00000018";
    when 16#2F3E# => romdata <= X"00000A98";
    when 16#2F3F# => romdata <= X"FFFFD6A4";
    when 16#2F40# => romdata <= X"00000104";
    when 16#2F41# => romdata <= X"00410D1E";
    when 16#2F42# => romdata <= X"2D45090F";
    when 16#2F43# => romdata <= X"1F000000";
    when 16#2F44# => romdata <= X"00000010";
    when 16#2F45# => romdata <= X"00000AB4";
    when 16#2F46# => romdata <= X"FFFFD78C";
    when 16#2F47# => romdata <= X"00000034";
    when 16#2F49# => romdata <= X"00000010";
    when 16#2F4A# => romdata <= X"00000AC8";
    when 16#2F4B# => romdata <= X"FFFFD7AC";
    when 16#2F4C# => romdata <= X"00000028";
    when 16#2F4E# => romdata <= X"00000010";
    when 16#2F4F# => romdata <= X"00000ADC";
    when 16#2F50# => romdata <= X"FFFFD7C0";
    when 16#2F51# => romdata <= X"0000001C";
    when 16#2F53# => romdata <= X"00000018";
    when 16#2F54# => romdata <= X"00000AF0";
    when 16#2F55# => romdata <= X"FFFFD7C8";
    when 16#2F56# => romdata <= X"00000058";
    when 16#2F57# => romdata <= X"00410D1E";
    when 16#2F58# => romdata <= X"2D44090F";
    when 16#2F59# => romdata <= X"1F000000";
    when 16#2F5A# => romdata <= X"00000018";
    when 16#2F5B# => romdata <= X"00000B0C";
    when 16#2F5C# => romdata <= X"FFFFD804";
    when 16#2F5D# => romdata <= X"00000058";
    when 16#2F5E# => romdata <= X"00410D1E";
    when 16#2F5F# => romdata <= X"2D4A090F";
    when 16#2F60# => romdata <= X"1F000000";
    when 16#2F61# => romdata <= X"00000018";
    when 16#2F62# => romdata <= X"00000B28";
    when 16#2F63# => romdata <= X"FFFFD840";
    when 16#2F64# => romdata <= X"00000050";
    when 16#2F65# => romdata <= X"00410D1E";
    when 16#2F66# => romdata <= X"2D44090F";
    when 16#2F67# => romdata <= X"1F000000";
    when 16#2F68# => romdata <= X"00000018";
    when 16#2F69# => romdata <= X"00000B44";
    when 16#2F6A# => romdata <= X"FFFFD874";
    when 16#2F6B# => romdata <= X"00000094";
    when 16#2F6C# => romdata <= X"00410D1E";
    when 16#2F6D# => romdata <= X"2D5D090F";
    when 16#2F6E# => romdata <= X"1F000000";
    when 16#2F6F# => romdata <= X"00000018";
    when 16#2F70# => romdata <= X"00000B60";
    when 16#2F71# => romdata <= X"FFFFD8EC";
    when 16#2F72# => romdata <= X"00000048";
    when 16#2F73# => romdata <= X"00410D1E";
    when 16#2F74# => romdata <= X"2D44090F";
    when 16#2F75# => romdata <= X"1F000000";
    when 16#2F76# => romdata <= X"00000018";
    when 16#2F77# => romdata <= X"00000B7C";
    when 16#2F78# => romdata <= X"FFFFD918";
    when 16#2F79# => romdata <= X"000000A0";
    when 16#2F7A# => romdata <= X"00410D1E";
    when 16#2F7B# => romdata <= X"2D41090F";
    when 16#2F7C# => romdata <= X"1F000000";
    when 16#2F7D# => romdata <= X"00000018";
    when 16#2F7E# => romdata <= X"00000B98";
    when 16#2F7F# => romdata <= X"FFFFD99C";
    when 16#2F80# => romdata <= X"00000040";
    when 16#2F81# => romdata <= X"00410D1E";
    when 16#2F82# => romdata <= X"2D42090F";
    when 16#2F83# => romdata <= X"1F000000";
    when 16#2F84# => romdata <= X"00000018";
    when 16#2F85# => romdata <= X"00000BB4";
    when 16#2F86# => romdata <= X"FFFFD9C0";
    when 16#2F87# => romdata <= X"00000170";
    when 16#2F88# => romdata <= X"00410D1E";
    when 16#2F89# => romdata <= X"2D43090F";
    when 16#2F8A# => romdata <= X"1F000000";
    when 16#2F8B# => romdata <= X"00000010";
    when 16#2F8C# => romdata <= X"00000BD0";
    when 16#2F8D# => romdata <= X"FFFFDB14";
    when 16#2F8E# => romdata <= X"0000001C";
    when 16#2F90# => romdata <= X"00000018";
    when 16#2F91# => romdata <= X"00000BE4";
    when 16#2F92# => romdata <= X"FFFFDB1C";
    when 16#2F93# => romdata <= X"00000044";
    when 16#2F94# => romdata <= X"00410D1E";
    when 16#2F95# => romdata <= X"2D43090F";
    when 16#2F96# => romdata <= X"1F000000";
    when 16#2F97# => romdata <= X"00000018";
    when 16#2F98# => romdata <= X"00000C00";
    when 16#2F99# => romdata <= X"FFFFDB44";
    when 16#2F9A# => romdata <= X"00000048";
    when 16#2F9B# => romdata <= X"00410D1E";
    when 16#2F9C# => romdata <= X"2D44090F";
    when 16#2F9D# => romdata <= X"1F000000";
    when 16#2F9E# => romdata <= X"00000018";
    when 16#2F9F# => romdata <= X"00000C1C";
    when 16#2FA0# => romdata <= X"FFFFDB70";
    when 16#2FA1# => romdata <= X"00000048";
    when 16#2FA2# => romdata <= X"00410D1E";
    when 16#2FA3# => romdata <= X"2D44090F";
    when 16#2FA4# => romdata <= X"1F000000";
    when 16#2FA5# => romdata <= X"00000010";
    when 16#2FA6# => romdata <= X"00000C38";
    when 16#2FA7# => romdata <= X"FFFFE1E4";
    when 16#2FA8# => romdata <= X"00000008";
    when 16#2FAA# => romdata <= X"00000010";
    when 16#2FAB# => romdata <= X"00000C4C";
    when 16#2FAC# => romdata <= X"FFFFE1D8";
    when 16#2FAD# => romdata <= X"00000014";
    when 16#2FAF# => romdata <= X"00000010";
    when 16#2FB0# => romdata <= X"00000C60";
    when 16#2FB1# => romdata <= X"FFFFE1D8";
    when 16#2FB2# => romdata <= X"00000008";
    when 16#2FB4# => romdata <= X"00000014";
    when 16#2FB5# => romdata <= X"00000C74";
    when 16#2FB6# => romdata <= X"FFFFE1CC";
    when 16#2FB7# => romdata <= X"0000001C";
    when 16#2FB8# => romdata <= X"00410D1E";
    when 16#2FB9# => romdata <= X"2D090F1F";
    when 16#2FBA# => romdata <= X"00000018";
    when 16#2FBB# => romdata <= X"00000C8C";
    when 16#2FBC# => romdata <= X"FFFFE1D0";
    when 16#2FBD# => romdata <= X"0000005C";
    when 16#2FBE# => romdata <= X"00410D1E";
    when 16#2FBF# => romdata <= X"2D44090F";
    when 16#2FC0# => romdata <= X"1F000000";
    when 16#2FC1# => romdata <= X"00000010";
    when 16#2FC2# => romdata <= X"00000CA8";
    when 16#2FC3# => romdata <= X"FFFFE210";
    when 16#2FC4# => romdata <= X"0000003C";
    when 16#2FC6# => romdata <= X"00000018";
    when 16#2FC7# => romdata <= X"00000CBC";
    when 16#2FC8# => romdata <= X"FFFFE238";
    when 16#2FC9# => romdata <= X"00000078";
    when 16#2FCA# => romdata <= X"00410D1E";
    when 16#2FCB# => romdata <= X"2D45090F";
    when 16#2FCC# => romdata <= X"1F000000";
    when 16#2FCD# => romdata <= X"00000010";
    when 16#2FCE# => romdata <= X"00000CD8";
    when 16#2FCF# => romdata <= X"FFFFE294";
    when 16#2FD0# => romdata <= X"00000050";
    when 16#2FD2# => romdata <= X"00000010";
    when 16#2FD3# => romdata <= X"00000CEC";
    when 16#2FD4# => romdata <= X"FFFFE2D0";
    when 16#2FD5# => romdata <= X"00000034";
    when 16#2FD7# => romdata <= X"00000018";
    when 16#2FD8# => romdata <= X"00000D00";
    when 16#2FD9# => romdata <= X"FFFFE7C0";
    when 16#2FDA# => romdata <= X"00000088";
    when 16#2FDB# => romdata <= X"00410D1E";
    when 16#2FDC# => romdata <= X"2D52090F";
    when 16#2FDD# => romdata <= X"1F000000";
    when 16#2FDE# => romdata <= X"00000010";
    when 16#2FDF# => romdata <= X"00000D1C";
    when 16#2FE0# => romdata <= X"FFFFE82C";
    when 16#2FE1# => romdata <= X"0000001C";
    when 16#2FE3# => romdata <= X"00000018";
    when 16#2FE4# => romdata <= X"00000D30";
    when 16#2FE5# => romdata <= X"FFFFE834";
    when 16#2FE6# => romdata <= X"00000120";
    when 16#2FE7# => romdata <= X"00410D1E";
    when 16#2FE8# => romdata <= X"2D58090F";
    when 16#2FE9# => romdata <= X"1F000000";
    when 16#2FEA# => romdata <= X"00000010";
    when 16#2FEB# => romdata <= X"00000D4C";
    when 16#2FEC# => romdata <= X"FFFFEA70";
    when 16#2FED# => romdata <= X"00000010";
    when 16#2FEF# => romdata <= X"00000018";
    when 16#2FF0# => romdata <= X"00000D60";
    when 16#2FF1# => romdata <= X"FFFFEA6C";
    when 16#2FF2# => romdata <= X"00000034";
    when 16#2FF3# => romdata <= X"00410D1E";
    when 16#2FF4# => romdata <= X"2D47090F";
    when 16#2FF5# => romdata <= X"1F000000";
    when 16#2FF6# => romdata <= X"00000018";
    when 16#2FF7# => romdata <= X"00000D7C";
    when 16#2FF8# => romdata <= X"FFFFEA84";
    when 16#2FF9# => romdata <= X"0000002C";
    when 16#2FFA# => romdata <= X"00410D1E";
    when 16#2FFB# => romdata <= X"2D45090F";
    when 16#2FFC# => romdata <= X"1F000000";
    when 16#2FFD# => romdata <= X"00000018";
    when 16#2FFE# => romdata <= X"00000D98";
    when 16#2FFF# => romdata <= X"FFFFEA94";
    when 16#3000# => romdata <= X"0000002C";
    when 16#3001# => romdata <= X"00410D1E";
    when 16#3002# => romdata <= X"2D45090F";
    when 16#3003# => romdata <= X"1F000000";
    when 16#3004# => romdata <= X"00000018";
    when 16#3005# => romdata <= X"00000DB4";
    when 16#3006# => romdata <= X"FFFFEAA4";
    when 16#3007# => romdata <= X"0000002C";
    when 16#3008# => romdata <= X"00410D1E";
    when 16#3009# => romdata <= X"2D45090F";
    when 16#300A# => romdata <= X"1F000000";
    when 16#300B# => romdata <= X"00000018";
    when 16#300C# => romdata <= X"00000DD0";
    when 16#300D# => romdata <= X"FFFFEAB4";
    when 16#300E# => romdata <= X"0000002C";
    when 16#300F# => romdata <= X"00410D1E";
    when 16#3010# => romdata <= X"2D45090F";
    when 16#3011# => romdata <= X"1F000000";
    when 16#3012# => romdata <= X"00000018";
    when 16#3013# => romdata <= X"00000DEC";
    when 16#3014# => romdata <= X"FFFFEAC4";
    when 16#3015# => romdata <= X"0000002C";
    when 16#3016# => romdata <= X"00410D1E";
    when 16#3017# => romdata <= X"2D45090F";
    when 16#3018# => romdata <= X"1F000000";
    when 16#3019# => romdata <= X"00000018";
    when 16#301A# => romdata <= X"00000E08";
    when 16#301B# => romdata <= X"FFFFEAD4";
    when 16#301C# => romdata <= X"0000002C";
    when 16#301D# => romdata <= X"00410D1E";
    when 16#301E# => romdata <= X"2D45090F";
    when 16#301F# => romdata <= X"1F000000";
    when 16#3020# => romdata <= X"00000018";
    when 16#3021# => romdata <= X"00000E24";
    when 16#3022# => romdata <= X"FFFFEAE4";
    when 16#3023# => romdata <= X"00000034";
    when 16#3024# => romdata <= X"00410D1E";
    when 16#3025# => romdata <= X"2D47090F";
    when 16#3026# => romdata <= X"1F000000";
    when 16#3027# => romdata <= X"00000018";
    when 16#3028# => romdata <= X"00000E40";
    when 16#3029# => romdata <= X"FFFFECA8";
    when 16#302A# => romdata <= X"0000004C";
    when 16#302B# => romdata <= X"00410D1E";
    when 16#302C# => romdata <= X"2D47090F";
    when 16#302D# => romdata <= X"1F000000";
    when 16#302E# => romdata <= X"00000010";
    when 16#302F# => romdata <= X"00000E5C";
    when 16#3030# => romdata <= X"FFFFF148";
    when 16#3031# => romdata <= X"0000000C";
    when 16#3034# => romdata <= X"00000004";
    when 16#3035# => romdata <= X"FFFFFFFF";
    when 16#3036# => romdata <= X"400023F8";
    when 16#3037# => romdata <= X"400024FC";
    when 16#303A# => romdata <= X"00000002";
    when 16#303B# => romdata <= X"FFFFFFFF";
    when 16#303E# => romdata <= X"474E5353";
    when 16#303F# => romdata <= X"20696E74";
    when 16#3040# => romdata <= X"65727275";
    when 16#3041# => romdata <= X"70742068";
    when 16#3042# => romdata <= X"616E646C";
    when 16#3043# => romdata <= X"65723A20";
    when 16#3044# => romdata <= X"25640D0A";
    when 16#3046# => romdata <= X"49525134";
    when 16#3047# => romdata <= X"3A204750";
    when 16#3048# => romdata <= X"54696D65";
    when 16#3049# => romdata <= X"722C2025";
    when 16#304A# => romdata <= X"690D0A00";
    when 16#304C# => romdata <= X"45786563";
    when 16#304D# => romdata <= X"7574696F";
    when 16#304E# => romdata <= X"6E206272";
    when 16#304F# => romdata <= X"65616B0D";
    when 16#3050# => romdata <= X"0A000000";
    when 16#3052# => romdata <= X"476F746F";
    when 16#3053# => romdata <= X"20524F4D";
    when 16#3054# => romdata <= X"0D0A0000";
    when 16#3056# => romdata <= X"5245424F";
    when 16#3057# => romdata <= X"4F540D0A";
    when 16#305A# => romdata <= X"4C6F6164";
    when 16#305B# => romdata <= X"696E6720";
    when 16#305C# => romdata <= X"2E2E2E0D";
    when 16#305D# => romdata <= X"0A3E0000";
    when 16#305E# => romdata <= X"2441434B";
    when 16#305F# => romdata <= X"24000000";
    when 16#3060# => romdata <= X"426F6F74";
    when 16#3061# => romdata <= X"20466C61";
    when 16#3062# => romdata <= X"67203D20";
    when 16#3063# => romdata <= X"30782530";
    when 16#3064# => romdata <= X"38780D0A";
    when 16#3066# => romdata <= X"0D0A0D0A";
    when 16#3067# => romdata <= X"0D0A0D0A";
    when 16#3068# => romdata <= X"0D0A0D0A";
    when 16#3069# => romdata <= X"0D0A0D0A";
    when 16#306A# => romdata <= X"09465047";
    when 16#306B# => romdata <= X"412F4153";
    when 16#306C# => romdata <= X"49432076";
    when 16#306D# => romdata <= X"616C6964";
    when 16#306E# => romdata <= X"6174696F";
    when 16#306F# => romdata <= X"6E206669";
    when 16#3070# => romdata <= X"726D7761";
    when 16#3071# => romdata <= X"72652076";
    when 16#3072# => romdata <= X"2E302E39";
    when 16#3073# => romdata <= X"202F3230";
    when 16#3074# => romdata <= X"31322E30";
    when 16#3075# => romdata <= X"312E3331";
    when 16#3076# => romdata <= X"2F0D0A0D";
    when 16#3077# => romdata <= X"0A000000";
    when 16#3078# => romdata <= X"53656C65";
    when 16#3079# => romdata <= X"63742074";
    when 16#307A# => romdata <= X"65737420";
    when 16#307B# => romdata <= X"28707265";
    when 16#307C# => romdata <= X"7373206B";
    when 16#307D# => romdata <= X"6579626F";
    when 16#307E# => romdata <= X"61726420";
    when 16#307F# => romdata <= X"62757474";
    when 16#3080# => romdata <= X"6F6E293A";
    when 16#3081# => romdata <= X"0D0A0000";
    when 16#3082# => romdata <= X"09312E20";
    when 16#3083# => romdata <= X"52656164";
    when 16#3084# => romdata <= X"20626F6F";
    when 16#3085# => romdata <= X"7420666C";
    when 16#3086# => romdata <= X"61670D0A";
    when 16#3088# => romdata <= X"09322E20";
    when 16#3089# => romdata <= X"52656164";
    when 16#308A# => romdata <= X"20737973";
    when 16#308B# => romdata <= X"74656D20";
    when 16#308C# => romdata <= X"706C7567";
    when 16#308D# => romdata <= X"276E2770";
    when 16#308E# => romdata <= X"6C617920";
    when 16#308F# => romdata <= X"696E666F";
    when 16#3090# => romdata <= X"726D6174";
    when 16#3091# => romdata <= X"696F6E0D";
    when 16#3092# => romdata <= X"0A000000";
    when 16#3094# => romdata <= X"09332E20";
    when 16#3095# => romdata <= X"47505469";
    when 16#3096# => romdata <= X"6D657220";
    when 16#3097# => romdata <= X"496E7465";
    when 16#3098# => romdata <= X"72727570";
    when 16#3099# => romdata <= X"74207075";
    when 16#309A# => romdata <= X"6C736520";
    when 16#309B# => romdata <= X"64657465";
    when 16#309C# => romdata <= X"6374696F";
    when 16#309D# => romdata <= X"6E0D0A00";
    when 16#309E# => romdata <= X"09342E20";
    when 16#309F# => romdata <= X"474E5353";
    when 16#30A0# => romdata <= X"20456E67";
    when 16#30A1# => romdata <= X"696E6520";
    when 16#30A2# => romdata <= X"496E7465";
    when 16#30A3# => romdata <= X"72727570";
    when 16#30A4# => romdata <= X"74207075";
    when 16#30A5# => romdata <= X"6C736520";
    when 16#30A6# => romdata <= X"64657465";
    when 16#30A7# => romdata <= X"6374696F";
    when 16#30A8# => romdata <= X"6E0D0A00";
    when 16#30AA# => romdata <= X"09352E20";
    when 16#30AB# => romdata <= X"52656164";
    when 16#30AC# => romdata <= X"20474E53";
    when 16#30AD# => romdata <= X"53206D65";
    when 16#30AE# => romdata <= X"6D6F7279";
    when 16#30AF# => romdata <= X"0D0A0000";
    when 16#30B0# => romdata <= X"09626F6F";
    when 16#30B1# => romdata <= X"742E2043";
    when 16#30B2# => romdata <= X"6865636B";
    when 16#30B3# => romdata <= X"20666972";
    when 16#30B4# => romdata <= X"6D776172";
    when 16#30B5# => romdata <= X"65206C6F";
    when 16#30B6# => romdata <= X"61646572";
    when 16#30B7# => romdata <= X"2066756E";
    when 16#30B8# => romdata <= X"6374696F";
    when 16#30B9# => romdata <= X"6E616C69";
    when 16#30BA# => romdata <= X"74790D0A";
    when 16#30BC# => romdata <= X"09612E20";
    when 16#30BD# => romdata <= X"52756E20";
    when 16#30BE# => romdata <= X"616C6C20";
    when 16#30BF# => romdata <= X"74657374";
    when 16#30C0# => romdata <= X"730D0A00";
    when 16#30C2# => romdata <= X"0D0A3E00";
    when 16#30C4# => romdata <= X"474E5353";
    when 16#30C5# => romdata <= X"20456E67";
    when 16#30C6# => romdata <= X"696E6520";
    when 16#30C7# => romdata <= X"6D656D6F";
    when 16#30C8# => romdata <= X"72793A0D";
    when 16#30C9# => romdata <= X"0A000000";
    when 16#30CA# => romdata <= X"5B253038";
    when 16#30CB# => romdata <= X"785D2030";
    when 16#30CC# => romdata <= X"78253038";
    when 16#30CD# => romdata <= X"780D0A00";
    when 16#30CE# => romdata <= X"4761696C";
    when 16#30CF# => romdata <= X"73657220";
    when 16#30D0# => romdata <= X"5648444C";
    when 16#30D1# => romdata <= X"206C6962";
    when 16#30D2# => romdata <= X"72617279";
    when 16#30D3# => romdata <= X"20627569";
    when 16#30D4# => romdata <= X"6C643A20";
    when 16#30D5# => romdata <= X"25640D0A";
    when 16#30D8# => romdata <= X"44657669";
    when 16#30D9# => romdata <= X"63652049";
    when 16#30DA# => romdata <= X"443A2030";
    when 16#30DB# => romdata <= X"78253034";
    when 16#30DC# => romdata <= X"780D0A0D";
    when 16#30DD# => romdata <= X"0A000000";
    when 16#30DE# => romdata <= X"25732009";
    when 16#30DF# => romdata <= X"09202725";
    when 16#30E0# => romdata <= X"73273A0D";
    when 16#30E1# => romdata <= X"0A000000";
    when 16#30E2# => romdata <= X"20202020";
    when 16#30E3# => romdata <= X"41484220";
    when 16#30E4# => romdata <= X"6D617374";
    when 16#30E5# => romdata <= X"65725B25";
    when 16#30E6# => romdata <= X"645D3A20";
    when 16#30E7# => romdata <= X"7665722E";
    when 16#30E8# => romdata <= X"2025690D";
    when 16#30E9# => romdata <= X"0A000000";
    when 16#30EA# => romdata <= X"20202020";
    when 16#30EB# => romdata <= X"736C765B";
    when 16#30EC# => romdata <= X"25645D3A";
    when 16#30ED# => romdata <= X"20307825";
    when 16#30EE# => romdata <= X"3038782E";
    when 16#30EF# => romdata <= X"2E307825";
    when 16#30F0# => romdata <= X"3038780D";
    when 16#30F1# => romdata <= X"0A000000";
    when 16#30F2# => romdata <= X"25732009";
    when 16#30F3# => romdata <= X"09202725";
    when 16#30F4# => romdata <= X"73270D0A";
    when 16#30F6# => romdata <= X"20202020";
    when 16#30F7# => romdata <= X"6170625B";
    when 16#30F8# => romdata <= X"25645D20";
    when 16#30F9# => romdata <= X"30782530";
    when 16#30FA# => romdata <= X"38782E2E";
    when 16#30FB# => romdata <= X"30782530";
    when 16#30FC# => romdata <= X"38780D0A";
    when 16#30FE# => romdata <= X"474E5353";
    when 16#30FF# => romdata <= X"20696E74";
    when 16#3100# => romdata <= X"65727275";
    when 16#3101# => romdata <= X"70742065";
    when 16#3102# => romdata <= X"6E61626C";
    when 16#3103# => romdata <= X"653A0D0A";
    when 16#3106# => romdata <= X"4E756D62";
    when 16#3107# => romdata <= X"6572206F";
    when 16#3108# => romdata <= X"6620696E";
    when 16#3109# => romdata <= X"74657272";
    when 16#310A# => romdata <= X"75707473";
    when 16#310B# => romdata <= X"3A202020";
    when 16#310C# => romdata <= X"25692F25";
    when 16#310D# => romdata <= X"690D0A00";
    when 16#310E# => romdata <= X"474E5353";
    when 16#310F# => romdata <= X"20696E74";
    when 16#3110# => romdata <= X"65727275";
    when 16#3111# => romdata <= X"70742064";
    when 16#3112# => romdata <= X"69736162";
    when 16#3113# => romdata <= X"6C652E0D";
    when 16#3114# => romdata <= X"0A000000";
    when 16#3116# => romdata <= X"47505469";
    when 16#3117# => romdata <= X"6D657220";
    when 16#3118# => romdata <= X"696E7465";
    when 16#3119# => romdata <= X"72727570";
    when 16#311A# => romdata <= X"7420656E";
    when 16#311B# => romdata <= X"61626C65";
    when 16#311C# => romdata <= X"3A0D0A00";
    when 16#311E# => romdata <= X"4E756D62";
    when 16#311F# => romdata <= X"6572206F";
    when 16#3120# => romdata <= X"6620696E";
    when 16#3121# => romdata <= X"74657272";
    when 16#3122# => romdata <= X"75707473";
    when 16#3123# => romdata <= X"3A202020";
    when 16#3124# => romdata <= X"25690D0A";
    when 16#3126# => romdata <= X"47505469";
    when 16#3127# => romdata <= X"6D657220";
    when 16#3128# => romdata <= X"696E7465";
    when 16#3129# => romdata <= X"72727570";
    when 16#312A# => romdata <= X"74206469";
    when 16#312B# => romdata <= X"7361626C";
    when 16#312C# => romdata <= X"653A0D0A";
    when 16#312E# => romdata <= X"31000000";
    when 16#3130# => romdata <= X"32000000";
    when 16#3132# => romdata <= X"33000000";
    when 16#3134# => romdata <= X"34000000";
    when 16#3136# => romdata <= X"35000000";
    when 16#3138# => romdata <= X"626F6F74";
    when 16#313A# => romdata <= X"61000000";
    when 16#313C# => romdata <= X"596F7520";
    when 16#313D# => romdata <= X"7072696E";
    when 16#313E# => romdata <= X"74202225";
    when 16#313F# => romdata <= X"73220D0A";
    when 16#3142# => romdata <= X"0D0A5072";
    when 16#3143# => romdata <= X"65737320";
    when 16#3144# => romdata <= X"27456E74";
    when 16#3145# => romdata <= X"65722720";
    when 16#3146# => romdata <= X"746F2063";
    when 16#3147# => romdata <= X"6F6E7469";
    when 16#3148# => romdata <= X"6E756520";
    when 16#3149# => romdata <= X"6F722027";
    when 16#314A# => romdata <= X"72272074";
    when 16#314B# => romdata <= X"6F207265";
    when 16#314C# => romdata <= X"70656164";
    when 16#314D# => romdata <= X"20746573";
    when 16#314E# => romdata <= X"74202E20";
    when 16#314F# => romdata <= X"2E202E0D";
    when 16#3150# => romdata <= X"0A3E0000";
    when 16#3152# => romdata <= X"556E6B6E";
    when 16#3153# => romdata <= X"6F776E20";
    when 16#3154# => romdata <= X"20202020";
    when 16#3155# => romdata <= X"20202020";
    when 16#3156# => romdata <= X"20202020";
    when 16#3157# => romdata <= X"20202020";
    when 16#3158# => romdata <= X"20202020";
    when 16#3159# => romdata <= X"20202000";
    when 16#315A# => romdata <= X"43505520";
    when 16#315B# => romdata <= X"4C656F6E";
    when 16#315C# => romdata <= X"33202020";
    when 16#315D# => romdata <= X"20202020";
    when 16#315E# => romdata <= X"20202020";
    when 16#315F# => romdata <= X"20202020";
    when 16#3160# => romdata <= X"20202020";
    when 16#3161# => romdata <= X"20202000";
    when 16#3162# => romdata <= X"4C454F4E";
    when 16#3163# => romdata <= X"33204465";
    when 16#3164# => romdata <= X"62756720";
    when 16#3165# => romdata <= X"53757070";
    when 16#3166# => romdata <= X"6F727420";
    when 16#3167# => romdata <= X"556E6974";
    when 16#3168# => romdata <= X"20202020";
    when 16#3169# => romdata <= X"20202000";
    when 16#316A# => romdata <= X"4148422F";
    when 16#316B# => romdata <= X"41504220";
    when 16#316C# => romdata <= X"62726964";
    when 16#316D# => romdata <= X"67652020";
    when 16#316E# => romdata <= X"20202020";
    when 16#316F# => romdata <= X"20202020";
    when 16#3170# => romdata <= X"20202020";
    when 16#3171# => romdata <= X"20202000";
    when 16#3172# => romdata <= X"41504220";
    when 16#3173# => romdata <= X"55415254";
    when 16#3174# => romdata <= X"20202020";
    when 16#3175# => romdata <= X"20202020";
    when 16#3176# => romdata <= X"20202020";
    when 16#3177# => romdata <= X"20202020";
    when 16#3178# => romdata <= X"20202020";
    when 16#3179# => romdata <= X"20202000";
    when 16#317A# => romdata <= X"4D756C74";
    when 16#317B# => romdata <= X"692D7072";
    when 16#317C# => romdata <= X"6F636573";
    when 16#317D# => romdata <= X"736F7220";
    when 16#317E# => romdata <= X"49525120";
    when 16#317F# => romdata <= X"636F6E74";
    when 16#3180# => romdata <= X"726F6C6C";
    when 16#3181# => romdata <= X"65722000";
    when 16#3182# => romdata <= X"41484220";
    when 16#3183# => romdata <= X"5352414D";
    when 16#3184# => romdata <= X"20202020";
    when 16#3185# => romdata <= X"20202020";
    when 16#3186# => romdata <= X"20202020";
    when 16#3187# => romdata <= X"20202020";
    when 16#3188# => romdata <= X"20202020";
    when 16#3189# => romdata <= X"20202000";
    when 16#318A# => romdata <= X"47656E65";
    when 16#318B# => romdata <= X"72616C20";
    when 16#318C# => romdata <= X"50757270";
    when 16#318D# => romdata <= X"6F736520";
    when 16#318E# => romdata <= X"54696D65";
    when 16#318F# => romdata <= X"72732020";
    when 16#3190# => romdata <= X"20202020";
    when 16#3191# => romdata <= X"20202000";
    when 16#3192# => romdata <= X"41484220";
    when 16#3193# => romdata <= X"524F4D20";
    when 16#3194# => romdata <= X"20202020";
    when 16#3195# => romdata <= X"20202020";
    when 16#3196# => romdata <= X"20202020";
    when 16#3197# => romdata <= X"20202020";
    when 16#3198# => romdata <= X"20202020";
    when 16#3199# => romdata <= X"20202000";
    when 16#319A# => romdata <= X"41484220";
    when 16#319B# => romdata <= X"4A544147";
    when 16#319C# => romdata <= X"20202020";
    when 16#319D# => romdata <= X"20202020";
    when 16#319E# => romdata <= X"20202020";
    when 16#319F# => romdata <= X"20202020";
    when 16#31A0# => romdata <= X"20202020";
    when 16#31A1# => romdata <= X"20202000";
    when 16#31A2# => romdata <= X"52462066";
    when 16#31A3# => romdata <= X"726F6E74";
    when 16#31A4# => romdata <= X"2D656E64";
    when 16#31A5# => romdata <= X"20636F6E";
    when 16#31A6# => romdata <= X"74726F6C";
    when 16#31A7# => romdata <= X"6C657220";
    when 16#31A8# => romdata <= X"20202020";
    when 16#31A9# => romdata <= X"20202000";
    when 16#31AA# => romdata <= X"474E5353";
    when 16#31AB# => romdata <= X"20456E67";
    when 16#31AC# => romdata <= X"696E6520";
    when 16#31AD# => romdata <= X"20202020";
    when 16#31AE# => romdata <= X"20202020";
    when 16#31AF# => romdata <= X"20202020";
    when 16#31B0# => romdata <= X"20202020";
    when 16#31B1# => romdata <= X"20202000";
    when 16#31B2# => romdata <= X"332D6178";
    when 16#31B3# => romdata <= X"69732047";
    when 16#31B4# => romdata <= X"79726F73";
    when 16#31B5# => romdata <= X"636F7065";
    when 16#31B6# => romdata <= X"20636F6E";
    when 16#31B7# => romdata <= X"74726F6C";
    when 16#31B8# => romdata <= X"6C657220";
    when 16#31B9# => romdata <= X"20202000";
    when 16#31BA# => romdata <= X"332D6178";
    when 16#31BB# => romdata <= X"69732041";
    when 16#31BC# => romdata <= X"6363656C";
    when 16#31BD# => romdata <= X"65726F6D";
    when 16#31BE# => romdata <= X"65746572";
    when 16#31BF# => romdata <= X"20636F6E";
    when 16#31C0# => romdata <= X"74726F6C";
    when 16#31C1# => romdata <= X"6C657200";
    when 16#31C2# => romdata <= X"4669726D";
    when 16#31C3# => romdata <= X"77617265";
    when 16#31C4# => romdata <= X"20524F4D";
    when 16#31C5# => romdata <= X"20696D61";
    when 16#31C6# => romdata <= X"67652020";
    when 16#31C7# => romdata <= X"20202020";
    when 16#31C8# => romdata <= X"20202020";
    when 16#31C9# => romdata <= X"20202000";
    when 16#31CA# => romdata <= X"556E6B6E";
    when 16#31CB# => romdata <= X"6F776E20";
    when 16#31CC# => romdata <= X"20202020";
    when 16#31CD# => romdata <= X"20202020";
    when 16#31D0# => romdata <= X"47616973";
    when 16#31D1# => romdata <= X"6C657220";
    when 16#31D2# => romdata <= X"52657365";
    when 16#31D3# => romdata <= X"61726368";
    when 16#31D6# => romdata <= X"474E5353";
    when 16#31D7# => romdata <= X"2053656E";
    when 16#31D8# => romdata <= X"736F7220";
    when 16#31D9# => romdata <= X"4C746420";
    when 16#31DC# => romdata <= X"4000C548";
    when 16#31DD# => romdata <= X"00000003";
    when 16#31DE# => romdata <= X"4000C568";
    when 16#31DF# => romdata <= X"00000004";
    when 16#31E0# => romdata <= X"4000C588";
    when 16#31E1# => romdata <= X"00000006";
    when 16#31E2# => romdata <= X"4000C5A8";
    when 16#31E3# => romdata <= X"0000000C";
    when 16#31E4# => romdata <= X"4000C5C8";
    when 16#31E5# => romdata <= X"0000000D";
    when 16#31E6# => romdata <= X"4000C5E8";
    when 16#31E7# => romdata <= X"0000000E";
    when 16#31E8# => romdata <= X"4000C608";
    when 16#31E9# => romdata <= X"00000011";
    when 16#31EA# => romdata <= X"4000C628";
    when 16#31EB# => romdata <= X"0000001B";
    when 16#31EC# => romdata <= X"4000C648";
    when 16#31ED# => romdata <= X"0000001C";
    when 16#31EE# => romdata <= X"4000C668";
    when 16#31EF# => romdata <= X"00000077";
    when 16#31F0# => romdata <= X"4000C688";
    when 16#31F1# => romdata <= X"00000078";
    when 16#31F2# => romdata <= X"4000C6A8";
    when 16#31F3# => romdata <= X"00000079";
    when 16#31F4# => romdata <= X"4000C6C8";
    when 16#31F5# => romdata <= X"0000007A";
    when 16#31F6# => romdata <= X"4000C6E8";
    when 16#31F7# => romdata <= X"0000007B";
    when 16#31F8# => romdata <= X"4000C708";
    when 16#31FA# => romdata <= X"4000C728";
    when 16#31FB# => romdata <= X"00000001";
    when 16#31FC# => romdata <= X"4000C740";
    when 16#31FD# => romdata <= X"000000F1";
    when 16#31FE# => romdata <= X"4000C758";
    when 16#31FF# => romdata <= X"4000CAD0";
    when 16#3200# => romdata <= X"43000000";
    when 16#3202# => romdata <= X"30313233";
    when 16#3203# => romdata <= X"34353637";
    when 16#3204# => romdata <= X"38394142";
    when 16#3205# => romdata <= X"43444546";
    when 16#3208# => romdata <= X"496E6600";
    when 16#320A# => romdata <= X"30313233";
    when 16#320B# => romdata <= X"34353637";
    when 16#320C# => romdata <= X"38396162";
    when 16#320D# => romdata <= X"63646566";
    when 16#3210# => romdata <= X"4E614E00";
    when 16#3212# => romdata <= X"30000000";
    when 16#3214# => romdata <= X"2E000000";
    when 16#3216# => romdata <= X"286E756C";
    when 16#3217# => romdata <= X"6C290000";
    when 16#321A# => romdata <= X"30303030";
    when 16#321B# => romdata <= X"30303030";
    when 16#321C# => romdata <= X"30303030";
    when 16#321D# => romdata <= X"30303030";
    when 16#321E# => romdata <= X"20202020";
    when 16#321F# => romdata <= X"20202020";
    when 16#3220# => romdata <= X"20202020";
    when 16#3221# => romdata <= X"20202020";
    when 16#3222# => romdata <= X"432D5554";
    when 16#3223# => romdata <= X"462D3800";
    when 16#3224# => romdata <= X"432D534A";
    when 16#3225# => romdata <= X"49530000";
    when 16#3226# => romdata <= X"432D4555";
    when 16#3227# => romdata <= X"434A5000";
    when 16#3228# => romdata <= X"432D4A49";
    when 16#3229# => romdata <= X"53000000";
    when 16#322A# => romdata <= X"496E6669";
    when 16#322B# => romdata <= X"6E697479";
    when 16#322E# => romdata <= X"41F00000";
    when 16#3230# => romdata <= X"3FF80000";
    when 16#3232# => romdata <= X"3FD287A7";
    when 16#3233# => romdata <= X"636F4361";
    when 16#3234# => romdata <= X"3FC68A28";
    when 16#3235# => romdata <= X"8B60C8B3";
    when 16#3236# => romdata <= X"3FD34413";
    when 16#3237# => romdata <= X"509F79FB";
    when 16#3238# => romdata <= X"3FF00000";
    when 16#323A# => romdata <= X"40240000";
    when 16#323C# => romdata <= X"401C0000";
    when 16#323E# => romdata <= X"40140000";
    when 16#3240# => romdata <= X"3FE00000";
    when 16#3242# => romdata <= X"49534F2D";
    when 16#3243# => romdata <= X"38383539";
    when 16#3244# => romdata <= X"2D310000";
    when 16#3246# => romdata <= X"4000C850";
    when 16#3247# => romdata <= X"4000C500";
    when 16#3248# => romdata <= X"4000C500";
    when 16#3249# => romdata <= X"4000C500";
    when 16#324A# => romdata <= X"4000C500";
    when 16#324B# => romdata <= X"4000C500";
    when 16#324C# => romdata <= X"4000C500";
    when 16#324D# => romdata <= X"4000C500";
    when 16#324E# => romdata <= X"4000C500";
    when 16#324F# => romdata <= X"4000C500";
    when 16#3250# => romdata <= X"7F7F7F7F";
    when 16#3251# => romdata <= X"7F7F7F7F";
    when 16#3252# => romdata <= X"4000C908";
    when 16#3254# => romdata <= X"3FF00000";
    when 16#3256# => romdata <= X"40240000";
    when 16#3258# => romdata <= X"40590000";
    when 16#325A# => romdata <= X"408F4000";
    when 16#325C# => romdata <= X"40C38800";
    when 16#325E# => romdata <= X"40F86A00";
    when 16#3260# => romdata <= X"412E8480";
    when 16#3262# => romdata <= X"416312D0";
    when 16#3264# => romdata <= X"4197D784";
    when 16#3266# => romdata <= X"41CDCD65";
    when 16#3268# => romdata <= X"4202A05F";
    when 16#3269# => romdata <= X"20000000";
    when 16#326A# => romdata <= X"42374876";
    when 16#326B# => romdata <= X"E8000000";
    when 16#326C# => romdata <= X"426D1A94";
    when 16#326D# => romdata <= X"A2000000";
    when 16#326E# => romdata <= X"42A2309C";
    when 16#326F# => romdata <= X"E5400000";
    when 16#3270# => romdata <= X"42D6BCC4";
    when 16#3271# => romdata <= X"1E900000";
    when 16#3272# => romdata <= X"430C6BF5";
    when 16#3273# => romdata <= X"26340000";
    when 16#3274# => romdata <= X"4341C379";
    when 16#3275# => romdata <= X"37E08000";
    when 16#3276# => romdata <= X"43763457";
    when 16#3277# => romdata <= X"85D8A000";
    when 16#3278# => romdata <= X"43ABC16D";
    when 16#3279# => romdata <= X"674EC800";
    when 16#327A# => romdata <= X"43E158E4";
    when 16#327B# => romdata <= X"60913D00";
    when 16#327C# => romdata <= X"4415AF1D";
    when 16#327D# => romdata <= X"78B58C40";
    when 16#327E# => romdata <= X"444B1AE4";
    when 16#327F# => romdata <= X"D6E2EF50";
    when 16#3280# => romdata <= X"4480F0CF";
    when 16#3281# => romdata <= X"064DD592";
    when 16#3282# => romdata <= X"44B52D02";
    when 16#3283# => romdata <= X"C7E14AF6";
    when 16#3284# => romdata <= X"44EA7843";
    when 16#3285# => romdata <= X"79D99DB4";
    when 16#3286# => romdata <= X"4341C379";
    when 16#3287# => romdata <= X"37E08000";
    when 16#3288# => romdata <= X"4693B8B5";
    when 16#3289# => romdata <= X"B5056E17";
    when 16#328A# => romdata <= X"4D384F03";
    when 16#328B# => romdata <= X"E93FF9F5";
    when 16#328C# => romdata <= X"5A827748";
    when 16#328D# => romdata <= X"F9301D32";
    when 16#328E# => romdata <= X"75154FDD";
    when 16#328F# => romdata <= X"7F73BF3C";
    when 16#3290# => romdata <= X"3C9CD2B2";
    when 16#3291# => romdata <= X"97D889BC";
    when 16#3292# => romdata <= X"3949F623";
    when 16#3293# => romdata <= X"D5A8A733";
    when 16#3294# => romdata <= X"32A50FFD";
    when 16#3295# => romdata <= X"44F4A73D";
    when 16#3296# => romdata <= X"255BBA08";
    when 16#3297# => romdata <= X"CF8C979D";
    when 16#3298# => romdata <= X"0AC80628";
    when 16#3299# => romdata <= X"64AC6F43";
    when 16#329A# => romdata <= X"00000005";
    when 16#329B# => romdata <= X"00000019";
    when 16#329C# => romdata <= X"0000007D";
    when 16#329E# => romdata <= X"9DE3BFA0";
    when 16#329F# => romdata <= X"7FFFD1AB";
    when 16#32A0# => romdata <= X"01000000";
    when 16#32A1# => romdata <= X"7FFFF9E4";
    when 16#32A2# => romdata <= X"01000000";
    when 16#32A3# => romdata <= X"81C7E008";
    when 16#32A4# => romdata <= X"81E80000";
    when 16#32A5# => romdata <= X"9DE3BFA0";
    when 16#32A6# => romdata <= X"7FFFD179";
    when 16#32A7# => romdata <= X"01000000";
    when 16#32A8# => romdata <= X"81C7E008";
    when 16#32A9# => romdata <= X"81E80000";
    when 16#32AC# => romdata <= X"00000001";
    when 16#32B0# => romdata <= X"4000D858";
    when 16#32B2# => romdata <= X"4000CAD0";
    when 16#32B5# => romdata <= X"4000CDBC";
    when 16#32B6# => romdata <= X"4000CE88";
    when 16#32B7# => romdata <= X"4000CF54";
    when 16#32C1# => romdata <= X"4000C800";
    when 16#32DF# => romdata <= X"00000001";
    when 16#32E0# => romdata <= X"330EABCD";
    when 16#32E1# => romdata <= X"1234E66D";
    when 16#32E2# => romdata <= X"DEEC0005";
    when 16#32E3# => romdata <= X"000B0000";
    when 16#340A# => romdata <= X"4000D020";
    when 16#340B# => romdata <= X"4000D020";
    when 16#340C# => romdata <= X"4000D028";
    when 16#340D# => romdata <= X"4000D028";
    when 16#340E# => romdata <= X"4000D030";
    when 16#340F# => romdata <= X"4000D030";
    when 16#3410# => romdata <= X"4000D038";
    when 16#3411# => romdata <= X"4000D038";
    when 16#3412# => romdata <= X"4000D040";
    when 16#3413# => romdata <= X"4000D040";
    when 16#3414# => romdata <= X"4000D048";
    when 16#3415# => romdata <= X"4000D048";
    when 16#3416# => romdata <= X"4000D050";
    when 16#3417# => romdata <= X"4000D050";
    when 16#3418# => romdata <= X"4000D058";
    when 16#3419# => romdata <= X"4000D058";
    when 16#341A# => romdata <= X"4000D060";
    when 16#341B# => romdata <= X"4000D060";
    when 16#341C# => romdata <= X"4000D068";
    when 16#341D# => romdata <= X"4000D068";
    when 16#341E# => romdata <= X"4000D070";
    when 16#341F# => romdata <= X"4000D070";
    when 16#3420# => romdata <= X"4000D078";
    when 16#3421# => romdata <= X"4000D078";
    when 16#3422# => romdata <= X"4000D080";
    when 16#3423# => romdata <= X"4000D080";
    when 16#3424# => romdata <= X"4000D088";
    when 16#3425# => romdata <= X"4000D088";
    when 16#3426# => romdata <= X"4000D090";
    when 16#3427# => romdata <= X"4000D090";
    when 16#3428# => romdata <= X"4000D098";
    when 16#3429# => romdata <= X"4000D098";
    when 16#342A# => romdata <= X"4000D0A0";
    when 16#342B# => romdata <= X"4000D0A0";
    when 16#342C# => romdata <= X"4000D0A8";
    when 16#342D# => romdata <= X"4000D0A8";
    when 16#342E# => romdata <= X"4000D0B0";
    when 16#342F# => romdata <= X"4000D0B0";
    when 16#3430# => romdata <= X"4000D0B8";
    when 16#3431# => romdata <= X"4000D0B8";
    when 16#3432# => romdata <= X"4000D0C0";
    when 16#3433# => romdata <= X"4000D0C0";
    when 16#3434# => romdata <= X"4000D0C8";
    when 16#3435# => romdata <= X"4000D0C8";
    when 16#3436# => romdata <= X"4000D0D0";
    when 16#3437# => romdata <= X"4000D0D0";
    when 16#3438# => romdata <= X"4000D0D8";
    when 16#3439# => romdata <= X"4000D0D8";
    when 16#343A# => romdata <= X"4000D0E0";
    when 16#343B# => romdata <= X"4000D0E0";
    when 16#343C# => romdata <= X"4000D0E8";
    when 16#343D# => romdata <= X"4000D0E8";
    when 16#343E# => romdata <= X"4000D0F0";
    when 16#343F# => romdata <= X"4000D0F0";
    when 16#3440# => romdata <= X"4000D0F8";
    when 16#3441# => romdata <= X"4000D0F8";
    when 16#3442# => romdata <= X"4000D100";
    when 16#3443# => romdata <= X"4000D100";
    when 16#3444# => romdata <= X"4000D108";
    when 16#3445# => romdata <= X"4000D108";
    when 16#3446# => romdata <= X"4000D110";
    when 16#3447# => romdata <= X"4000D110";
    when 16#3448# => romdata <= X"4000D118";
    when 16#3449# => romdata <= X"4000D118";
    when 16#344A# => romdata <= X"4000D120";
    when 16#344B# => romdata <= X"4000D120";
    when 16#344C# => romdata <= X"4000D128";
    when 16#344D# => romdata <= X"4000D128";
    when 16#344E# => romdata <= X"4000D130";
    when 16#344F# => romdata <= X"4000D130";
    when 16#3450# => romdata <= X"4000D138";
    when 16#3451# => romdata <= X"4000D138";
    when 16#3452# => romdata <= X"4000D140";
    when 16#3453# => romdata <= X"4000D140";
    when 16#3454# => romdata <= X"4000D148";
    when 16#3455# => romdata <= X"4000D148";
    when 16#3456# => romdata <= X"4000D150";
    when 16#3457# => romdata <= X"4000D150";
    when 16#3458# => romdata <= X"4000D158";
    when 16#3459# => romdata <= X"4000D158";
    when 16#345A# => romdata <= X"4000D160";
    when 16#345B# => romdata <= X"4000D160";
    when 16#345C# => romdata <= X"4000D168";
    when 16#345D# => romdata <= X"4000D168";
    when 16#345E# => romdata <= X"4000D170";
    when 16#345F# => romdata <= X"4000D170";
    when 16#3460# => romdata <= X"4000D178";
    when 16#3461# => romdata <= X"4000D178";
    when 16#3462# => romdata <= X"4000D180";
    when 16#3463# => romdata <= X"4000D180";
    when 16#3464# => romdata <= X"4000D188";
    when 16#3465# => romdata <= X"4000D188";
    when 16#3466# => romdata <= X"4000D190";
    when 16#3467# => romdata <= X"4000D190";
    when 16#3468# => romdata <= X"4000D198";
    when 16#3469# => romdata <= X"4000D198";
    when 16#346A# => romdata <= X"4000D1A0";
    when 16#346B# => romdata <= X"4000D1A0";
    when 16#346C# => romdata <= X"4000D1A8";
    when 16#346D# => romdata <= X"4000D1A8";
    when 16#346E# => romdata <= X"4000D1B0";
    when 16#346F# => romdata <= X"4000D1B0";
    when 16#3470# => romdata <= X"4000D1B8";
    when 16#3471# => romdata <= X"4000D1B8";
    when 16#3472# => romdata <= X"4000D1C0";
    when 16#3473# => romdata <= X"4000D1C0";
    when 16#3474# => romdata <= X"4000D1C8";
    when 16#3475# => romdata <= X"4000D1C8";
    when 16#3476# => romdata <= X"4000D1D0";
    when 16#3477# => romdata <= X"4000D1D0";
    when 16#3478# => romdata <= X"4000D1D8";
    when 16#3479# => romdata <= X"4000D1D8";
    when 16#347A# => romdata <= X"4000D1E0";
    when 16#347B# => romdata <= X"4000D1E0";
    when 16#347C# => romdata <= X"4000D1E8";
    when 16#347D# => romdata <= X"4000D1E8";
    when 16#347E# => romdata <= X"4000D1F0";
    when 16#347F# => romdata <= X"4000D1F0";
    when 16#3480# => romdata <= X"4000D1F8";
    when 16#3481# => romdata <= X"4000D1F8";
    when 16#3482# => romdata <= X"4000D200";
    when 16#3483# => romdata <= X"4000D200";
    when 16#3484# => romdata <= X"4000D208";
    when 16#3485# => romdata <= X"4000D208";
    when 16#3486# => romdata <= X"4000D210";
    when 16#3487# => romdata <= X"4000D210";
    when 16#3488# => romdata <= X"4000D218";
    when 16#3489# => romdata <= X"4000D218";
    when 16#348A# => romdata <= X"4000D220";
    when 16#348B# => romdata <= X"4000D220";
    when 16#348C# => romdata <= X"4000D228";
    when 16#348D# => romdata <= X"4000D228";
    when 16#348E# => romdata <= X"4000D230";
    when 16#348F# => romdata <= X"4000D230";
    when 16#3490# => romdata <= X"4000D238";
    when 16#3491# => romdata <= X"4000D238";
    when 16#3492# => romdata <= X"4000D240";
    when 16#3493# => romdata <= X"4000D240";
    when 16#3494# => romdata <= X"4000D248";
    when 16#3495# => romdata <= X"4000D248";
    when 16#3496# => romdata <= X"4000D250";
    when 16#3497# => romdata <= X"4000D250";
    when 16#3498# => romdata <= X"4000D258";
    when 16#3499# => romdata <= X"4000D258";
    when 16#349A# => romdata <= X"4000D260";
    when 16#349B# => romdata <= X"4000D260";
    when 16#349C# => romdata <= X"4000D268";
    when 16#349D# => romdata <= X"4000D268";
    when 16#349E# => romdata <= X"4000D270";
    when 16#349F# => romdata <= X"4000D270";
    when 16#34A0# => romdata <= X"4000D278";
    when 16#34A1# => romdata <= X"4000D278";
    when 16#34A2# => romdata <= X"4000D280";
    when 16#34A3# => romdata <= X"4000D280";
    when 16#34A4# => romdata <= X"4000D288";
    when 16#34A5# => romdata <= X"4000D288";
    when 16#34A6# => romdata <= X"4000D290";
    when 16#34A7# => romdata <= X"4000D290";
    when 16#34A8# => romdata <= X"4000D298";
    when 16#34A9# => romdata <= X"4000D298";
    when 16#34AA# => romdata <= X"4000D2A0";
    when 16#34AB# => romdata <= X"4000D2A0";
    when 16#34AC# => romdata <= X"4000D2A8";
    when 16#34AD# => romdata <= X"4000D2A8";
    when 16#34AE# => romdata <= X"4000D2B0";
    when 16#34AF# => romdata <= X"4000D2B0";
    when 16#34B0# => romdata <= X"4000D2B8";
    when 16#34B1# => romdata <= X"4000D2B8";
    when 16#34B2# => romdata <= X"4000D2C0";
    when 16#34B3# => romdata <= X"4000D2C0";
    when 16#34B4# => romdata <= X"4000D2C8";
    when 16#34B5# => romdata <= X"4000D2C8";
    when 16#34B6# => romdata <= X"4000D2D0";
    when 16#34B7# => romdata <= X"4000D2D0";
    when 16#34B8# => romdata <= X"4000D2D8";
    when 16#34B9# => romdata <= X"4000D2D8";
    when 16#34BA# => romdata <= X"4000D2E0";
    when 16#34BB# => romdata <= X"4000D2E0";
    when 16#34BC# => romdata <= X"4000D2E8";
    when 16#34BD# => romdata <= X"4000D2E8";
    when 16#34BE# => romdata <= X"4000D2F0";
    when 16#34BF# => romdata <= X"4000D2F0";
    when 16#34C0# => romdata <= X"4000D2F8";
    when 16#34C1# => romdata <= X"4000D2F8";
    when 16#34C2# => romdata <= X"4000D300";
    when 16#34C3# => romdata <= X"4000D300";
    when 16#34C4# => romdata <= X"4000D308";
    when 16#34C5# => romdata <= X"4000D308";
    when 16#34C6# => romdata <= X"4000D310";
    when 16#34C7# => romdata <= X"4000D310";
    when 16#34C8# => romdata <= X"4000D318";
    when 16#34C9# => romdata <= X"4000D318";
    when 16#34CA# => romdata <= X"4000D320";
    when 16#34CB# => romdata <= X"4000D320";
    when 16#34CC# => romdata <= X"4000D328";
    when 16#34CD# => romdata <= X"4000D328";
    when 16#34CE# => romdata <= X"4000D330";
    when 16#34CF# => romdata <= X"4000D330";
    when 16#34D0# => romdata <= X"4000D338";
    when 16#34D1# => romdata <= X"4000D338";
    when 16#34D2# => romdata <= X"4000D340";
    when 16#34D3# => romdata <= X"4000D340";
    when 16#34D4# => romdata <= X"4000D348";
    when 16#34D5# => romdata <= X"4000D348";
    when 16#34D6# => romdata <= X"4000D350";
    when 16#34D7# => romdata <= X"4000D350";
    when 16#34D8# => romdata <= X"4000D358";
    when 16#34D9# => romdata <= X"4000D358";
    when 16#34DA# => romdata <= X"4000D360";
    when 16#34DB# => romdata <= X"4000D360";
    when 16#34DC# => romdata <= X"4000D368";
    when 16#34DD# => romdata <= X"4000D368";
    when 16#34DE# => romdata <= X"4000D370";
    when 16#34DF# => romdata <= X"4000D370";
    when 16#34E0# => romdata <= X"4000D378";
    when 16#34E1# => romdata <= X"4000D378";
    when 16#34E2# => romdata <= X"4000D380";
    when 16#34E3# => romdata <= X"4000D380";
    when 16#34E4# => romdata <= X"4000D388";
    when 16#34E5# => romdata <= X"4000D388";
    when 16#34E6# => romdata <= X"4000D390";
    when 16#34E7# => romdata <= X"4000D390";
    when 16#34E8# => romdata <= X"4000D398";
    when 16#34E9# => romdata <= X"4000D398";
    when 16#34EA# => romdata <= X"4000D3A0";
    when 16#34EB# => romdata <= X"4000D3A0";
    when 16#34EC# => romdata <= X"4000D3A8";
    when 16#34ED# => romdata <= X"4000D3A8";
    when 16#34EE# => romdata <= X"4000D3B0";
    when 16#34EF# => romdata <= X"4000D3B0";
    when 16#34F0# => romdata <= X"4000D3B8";
    when 16#34F1# => romdata <= X"4000D3B8";
    when 16#34F2# => romdata <= X"4000D3C0";
    when 16#34F3# => romdata <= X"4000D3C0";
    when 16#34F4# => romdata <= X"4000D3C8";
    when 16#34F5# => romdata <= X"4000D3C8";
    when 16#34F6# => romdata <= X"4000D3D0";
    when 16#34F7# => romdata <= X"4000D3D0";
    when 16#34F8# => romdata <= X"4000D3D8";
    when 16#34F9# => romdata <= X"4000D3D8";
    when 16#34FA# => romdata <= X"4000D3E0";
    when 16#34FB# => romdata <= X"4000D3E0";
    when 16#34FC# => romdata <= X"4000D3E8";
    when 16#34FD# => romdata <= X"4000D3E8";
    when 16#34FE# => romdata <= X"4000D3F0";
    when 16#34FF# => romdata <= X"4000D3F0";
    when 16#3500# => romdata <= X"4000D3F8";
    when 16#3501# => romdata <= X"4000D3F8";
    when 16#3502# => romdata <= X"4000D400";
    when 16#3503# => romdata <= X"4000D400";
    when 16#3504# => romdata <= X"4000D408";
    when 16#3505# => romdata <= X"4000D408";
    when 16#3506# => romdata <= X"4000D410";
    when 16#3507# => romdata <= X"4000D410";
    when 16#3508# => romdata <= X"4000D418";
    when 16#3509# => romdata <= X"4000D418";
    when 16#350A# => romdata <= X"00020000";
    when 16#350B# => romdata <= X"FFFFFFFF";
    when 16#350D# => romdata <= X"4000D430";
    when 16#3511# => romdata <= X"00000002";
    when 16#352A# => romdata <= X"4000D4A4";
    when 16#352E# => romdata <= X"00000002";
    when 16#3546# => romdata <= X"00000001";
    when 16#3548# => romdata <= X"43000000";
    when 16#357C# => romdata <= X"4000D550";
    when 16#357D# => romdata <= X"4000D550";
    when 16#3583# => romdata <= X"80000100";
    when 16#3584# => romdata <= X"00000008";
    when 16#3585# => romdata <= X"00000007";
    when 16#3586# => romdata <= X"00000006";
    when 16#3587# => romdata <= X"00000003";
    when 16#3589# => romdata <= X"FFFF8AD0";
    when 16#358A# => romdata <= X"80000310";
    when others => romdata <= (others => '0');
    end case;
  end process;
end;
